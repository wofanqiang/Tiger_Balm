module xpb_lut
(
    input logic [5:0] flag[57],
    output logic [255:0] xpb[57]
);
        
        
    always_comb begin
        case(flag[0])
            6'd0: xpb[0] = 256'd0;
            6'd1: xpb[0] = 256'd26959946667150639794667015087019630673716372585036390074623444647937;
            6'd2: xpb[0] = 256'd53919893334301279589334030174039261347432745170072780149246889295874;
            6'd3: xpb[0] = 256'd80879840001451919384001045261058892021149117755109170223870333943811;
            6'd4: xpb[0] = 256'd107839786668602559178668060348078522694865490340145560298493778591748;
            6'd5: xpb[0] = 256'd134799733335753198973335075435098153368581862925181950373117223239685;
            6'd6: xpb[0] = 256'd161759680002903838768002090522117784042298235510218340447740667887622;
            6'd7: xpb[0] = 256'd188719626670054478562669105609137414716014608095254730522364112535559;
            6'd8: xpb[0] = 256'd215679573337205118357336120696157045389730980680291120596987557183496;
            6'd9: xpb[0] = 256'd242639520004355758152003135783176676063447353265327510671611001831433;
            6'd10: xpb[0] = 256'd269599466671506397946670150870196306737163725850363900746234446479370;
            6'd11: xpb[0] = 256'd296559413338657037741337165957215937410880098435400290820857891127307;
            6'd12: xpb[0] = 256'd323519360005807677536004181044235568084596471020436680895481335775244;
            6'd13: xpb[0] = 256'd350479306672958317330671196131255198758312843605473070970104780423181;
            6'd14: xpb[0] = 256'd377439253340108957125338211218274829432029216190509461044728225071118;
            6'd15: xpb[0] = 256'd404399200007259596920005226305294460105745588775545851119351669719055;
            6'd16: xpb[0] = 256'd431359146674410236714672241392314090779461961360582241193975114366992;
            6'd17: xpb[0] = 256'd458319093341560876509339256479333721453178333945618631268598559014929;
            6'd18: xpb[0] = 256'd485279040008711516304006271566353352126894706530655021343222003662866;
            6'd19: xpb[0] = 256'd512238986675862156098673286653372982800611079115691411417845448310803;
            6'd20: xpb[0] = 256'd539198933343012795893340301740392613474327451700727801492468892958740;
            6'd21: xpb[0] = 256'd566158880010163435688007316827412244148043824285764191567092337606677;
            6'd22: xpb[0] = 256'd593118826677314075482674331914431874821760196870800581641715782254614;
            6'd23: xpb[0] = 256'd620078773344464715277341347001451505495476569455836971716339226902551;
            6'd24: xpb[0] = 256'd647038720011615355072008362088471136169192942040873361790962671550488;
            6'd25: xpb[0] = 256'd673998666678765994866675377175490766842909314625909751865586116198425;
            6'd26: xpb[0] = 256'd700958613345916634661342392262510397516625687210946141940209560846362;
            6'd27: xpb[0] = 256'd727918560013067274456009407349530028190342059795982532014833005494299;
            6'd28: xpb[0] = 256'd754878506680217914250676422436549658864058432381018922089456450142236;
            6'd29: xpb[0] = 256'd781838453347368554045343437523569289537774804966055312164079894790173;
            6'd30: xpb[0] = 256'd808798400014519193840010452610588920211491177551091702238703339438110;
            6'd31: xpb[0] = 256'd835758346681669833634677467697608550885207550136128092313326784086047;
            6'd32: xpb[0] = 256'd862718293348820473429344482784628181558923922721164482387950228733984;
            6'd33: xpb[0] = 256'd889678240015971113224011497871647812232640295306200872462573673381921;
            6'd34: xpb[0] = 256'd916638186683121753018678512958667442906356667891237262537197118029858;
            6'd35: xpb[0] = 256'd943598133350272392813345528045687073580073040476273652611820562677795;
            6'd36: xpb[0] = 256'd970558080017423032608012543132706704253789413061310042686444007325732;
            6'd37: xpb[0] = 256'd997518026684573672402679558219726334927505785646346432761067451973669;
            6'd38: xpb[0] = 256'd1024477973351724312197346573306745965601222158231382822835690896621606;
            6'd39: xpb[0] = 256'd1051437920018874951992013588393765596274938530816419212910314341269543;
            6'd40: xpb[0] = 256'd1078397866686025591786680603480785226948654903401455602984937785917480;
            6'd41: xpb[0] = 256'd1105357813353176231581347618567804857622371275986491993059561230565417;
            6'd42: xpb[0] = 256'd1132317760020326871376014633654824488296087648571528383134184675213354;
            6'd43: xpb[0] = 256'd1159277706687477511170681648741844118969804021156564773208808119861291;
            6'd44: xpb[0] = 256'd1186237653354628150965348663828863749643520393741601163283431564509228;
            6'd45: xpb[0] = 256'd1213197600021778790760015678915883380317236766326637553358055009157165;
            6'd46: xpb[0] = 256'd1240157546688929430554682694002903010990953138911673943432678453805102;
            6'd47: xpb[0] = 256'd1267117493356080070349349709089922641664669511496710333507301898453039;
            6'd48: xpb[0] = 256'd1294077440023230710144016724176942272338385884081746723581925343100976;
            6'd49: xpb[0] = 256'd1321037386690381349938683739263961903012102256666783113656548787748913;
            6'd50: xpb[0] = 256'd1347997333357531989733350754350981533685818629251819503731172232396850;
            6'd51: xpb[0] = 256'd1374957280024682629528017769438001164359535001836855893805795677044787;
            6'd52: xpb[0] = 256'd1401917226691833269322684784525020795033251374421892283880419121692724;
            6'd53: xpb[0] = 256'd1428877173358983909117351799612040425706967747006928673955042566340661;
            6'd54: xpb[0] = 256'd1455837120026134548912018814699060056380684119591965064029666010988598;
            6'd55: xpb[0] = 256'd1482797066693285188706685829786079687054400492177001454104289455636535;
            6'd56: xpb[0] = 256'd1509757013360435828501352844873099317728116864762037844178912900284472;
            6'd57: xpb[0] = 256'd1536716960027586468296019859960118948401833237347074234253536344932409;
            6'd58: xpb[0] = 256'd1563676906694737108090686875047138579075549609932110624328159789580346;
            6'd59: xpb[0] = 256'd1590636853361887747885353890134158209749265982517147014402783234228283;
            6'd60: xpb[0] = 256'd1617596800029038387680020905221177840422982355102183404477406678876220;
            6'd61: xpb[0] = 256'd1644556746696189027474687920308197471096698727687219794552030123524157;
            6'd62: xpb[0] = 256'd1671516693363339667269354935395217101770415100272256184626653568172094;
            6'd63: xpb[0] = 256'd1698476640030490307064021950482236732444131472857292574701277012820031;
        endcase
    end

    always_comb begin
        case(flag[1])
            6'd0: xpb[1] = 256'd0;
            6'd1: xpb[1] = 256'd1725436586697640946858688965569256363117847845442328964775900457467968;
            6'd2: xpb[1] = 256'd3450873173395281893717377931138512726235695690884657929551800914935936;
            6'd3: xpb[1] = 256'd5176309760092922840576066896707769089353543536326986894327701372403904;
            6'd4: xpb[1] = 256'd6901746346790563787434755862277025452471391381769315859103601829871872;
            6'd5: xpb[1] = 256'd8627182933488204734293444827846281815589239227211644823879502287339840;
            6'd6: xpb[1] = 256'd10352619520185845681152133793415538178707087072653973788655402744807808;
            6'd7: xpb[1] = 256'd12078056106883486628010822758984794541824934918096302753431303202275776;
            6'd8: xpb[1] = 256'd13803492693581127574869511724554050904942782763538631718207203659743744;
            6'd9: xpb[1] = 256'd15528929280278768521728200690123307268060630608980960682983104117211712;
            6'd10: xpb[1] = 256'd17254365866976409468586889655692563631178478454423289647759004574679680;
            6'd11: xpb[1] = 256'd18979802453674050415445578621261819994296326299865618612534905032147648;
            6'd12: xpb[1] = 256'd20705239040371691362304267586831076357414174145307947577310805489615616;
            6'd13: xpb[1] = 256'd22430675627069332309162956552400332720532021990750276542086705947083584;
            6'd14: xpb[1] = 256'd24156112213766973256021645517969589083649869836192605506862606404551552;
            6'd15: xpb[1] = 256'd25881548800464614202880334483538845446767717681634934471638506862019520;
            6'd16: xpb[1] = 256'd27606985387162255149739023449108101809885565527077263436414407319487488;
            6'd17: xpb[1] = 256'd29332421973859896096597712414677358173003413372519592401190307776955456;
            6'd18: xpb[1] = 256'd31057858560557537043456401380246614536121261217961921365966208234423424;
            6'd19: xpb[1] = 256'd32783295147255177990315090345815870899239109063404250330742108691891392;
            6'd20: xpb[1] = 256'd34508731733952818937173779311385127262356956908846579295518009149359360;
            6'd21: xpb[1] = 256'd36234168320650459884032468276954383625474804754288908260293909606827328;
            6'd22: xpb[1] = 256'd37959604907348100830891157242523639988592652599731237225069810064295296;
            6'd23: xpb[1] = 256'd39685041494045741777749846208092896351710500445173566189845710521763264;
            6'd24: xpb[1] = 256'd41410478080743382724608535173662152714828348290615895154621610979231232;
            6'd25: xpb[1] = 256'd43135914667441023671467224139231409077946196136058224119397511436699200;
            6'd26: xpb[1] = 256'd44861351254138664618325913104800665441064043981500553084173411894167168;
            6'd27: xpb[1] = 256'd46586787840836305565184602070369921804181891826942882048949312351635136;
            6'd28: xpb[1] = 256'd48312224427533946512043291035939178167299739672385211013725212809103104;
            6'd29: xpb[1] = 256'd50037661014231587458901980001508434530417587517827539978501113266571072;
            6'd30: xpb[1] = 256'd51763097600929228405760668967077690893535435363269868943277013724039040;
            6'd31: xpb[1] = 256'd53488534187626869352619357932646947256653283208712197908052914181507008;
            6'd32: xpb[1] = 256'd55213970774324510299478046898216203619771131054154526872828814638974976;
            6'd33: xpb[1] = 256'd56939407361022151246336735863785459982888978899596855837604715096442944;
            6'd34: xpb[1] = 256'd58664843947719792193195424829354716346006826745039184802380615553910912;
            6'd35: xpb[1] = 256'd60390280534417433140054113794923972709124674590481513767156516011378880;
            6'd36: xpb[1] = 256'd62115717121115074086912802760493229072242522435923842731932416468846848;
            6'd37: xpb[1] = 256'd63841153707812715033771491726062485435360370281366171696708316926314816;
            6'd38: xpb[1] = 256'd65566590294510355980630180691631741798478218126808500661484217383782784;
            6'd39: xpb[1] = 256'd67292026881207996927488869657200998161596065972250829626260117841250752;
            6'd40: xpb[1] = 256'd69017463467905637874347558622770254524713913817693158591036018298718720;
            6'd41: xpb[1] = 256'd70742900054603278821206247588339510887831761663135487555811918756186688;
            6'd42: xpb[1] = 256'd72468336641300919768064936553908767250949609508577816520587819213654656;
            6'd43: xpb[1] = 256'd74193773227998560714923625519478023614067457354020145485363719671122624;
            6'd44: xpb[1] = 256'd75919209814696201661782314485047279977185305199462474450139620128590592;
            6'd45: xpb[1] = 256'd77644646401393842608641003450616536340303153044904803414915520586058560;
            6'd46: xpb[1] = 256'd79370082988091483555499692416185792703421000890347132379691421043526528;
            6'd47: xpb[1] = 256'd81095519574789124502358381381755049066538848735789461344467321500994496;
            6'd48: xpb[1] = 256'd82820956161486765449217070347324305429656696581231790309243221958462464;
            6'd49: xpb[1] = 256'd84546392748184406396075759312893561792774544426674119274019122415930432;
            6'd50: xpb[1] = 256'd86271829334882047342934448278462818155892392272116448238795022873398400;
            6'd51: xpb[1] = 256'd87997265921579688289793137244032074519010240117558777203570923330866368;
            6'd52: xpb[1] = 256'd89722702508277329236651826209601330882128087963001106168346823788334336;
            6'd53: xpb[1] = 256'd91448139094974970183510515175170587245245935808443435133122724245802304;
            6'd54: xpb[1] = 256'd93173575681672611130369204140739843608363783653885764097898624703270272;
            6'd55: xpb[1] = 256'd94899012268370252077227893106309099971481631499328093062674525160738240;
            6'd56: xpb[1] = 256'd96624448855067893024086582071878356334599479344770422027450425618206208;
            6'd57: xpb[1] = 256'd98349885441765533970945271037447612697717327190212750992226326075674176;
            6'd58: xpb[1] = 256'd100075322028463174917803960003016869060835175035655079957002226533142144;
            6'd59: xpb[1] = 256'd101800758615160815864662648968586125423953022881097408921778126990610112;
            6'd60: xpb[1] = 256'd103526195201858456811521337934155381787070870726539737886554027448078080;
            6'd61: xpb[1] = 256'd105251631788556097758380026899724638150188718571982066851329927905546048;
            6'd62: xpb[1] = 256'd106977068375253738705238715865293894513306566417424395816105828363014016;
            6'd63: xpb[1] = 256'd108702504961951379652097404830863150876424414262866724780881728820481984;
        endcase
    end

    always_comb begin
        case(flag[2])
            6'd0: xpb[2] = 256'd0;
            6'd1: xpb[2] = 256'd110427941548649020598956093796432407239542262108309053745657629277949952;
            6'd2: xpb[2] = 256'd220855883097298041197912187592864814479084524216618107491315258555899904;
            6'd3: xpb[2] = 256'd331283824645947061796868281389297221718626786324927161236972887833849856;
            6'd4: xpb[2] = 256'd441711766194596082395824375185729628958169048433236214982630517111799808;
            6'd5: xpb[2] = 256'd552139707743245102994780468982162036197711310541545268728288146389749760;
            6'd6: xpb[2] = 256'd662567649291894123593736562778594443437253572649854322473945775667699712;
            6'd7: xpb[2] = 256'd772995590840543144192692656575026850676795834758163376219603404945649664;
            6'd8: xpb[2] = 256'd883423532389192164791648750371459257916338096866472429965261034223599616;
            6'd9: xpb[2] = 256'd993851473937841185390604844167891665155880358974781483710918663501549568;
            6'd10: xpb[2] = 256'd1104279415486490205989560937964324072395422621083090537456576292779499520;
            6'd11: xpb[2] = 256'd1214707357035139226588517031760756479634964883191399591202233922057449472;
            6'd12: xpb[2] = 256'd1325135298583788247187473125557188886874507145299708644947891551335399424;
            6'd13: xpb[2] = 256'd1435563240132437267786429219353621294114049407408017698693549180613349376;
            6'd14: xpb[2] = 256'd1545991181681086288385385313150053701353591669516326752439206809891299328;
            6'd15: xpb[2] = 256'd1656419123229735308984341406946486108593133931624635806184864439169249280;
            6'd16: xpb[2] = 256'd1766847064778384329583297500742918515832676193732944859930522068447199232;
            6'd17: xpb[2] = 256'd1877275006327033350182253594539350923072218455841253913676179697725149184;
            6'd18: xpb[2] = 256'd1987702947875682370781209688335783330311760717949562967421837327003099136;
            6'd19: xpb[2] = 256'd2098130889424331391380165782132215737551302980057872021167494956281049088;
            6'd20: xpb[2] = 256'd2208558830972980411979121875928648144790845242166181074913152585558999040;
            6'd21: xpb[2] = 256'd2318986772521629432578077969725080552030387504274490128658810214836948992;
            6'd22: xpb[2] = 256'd2429414714070278453177034063521512959269929766382799182404467844114898944;
            6'd23: xpb[2] = 256'd2539842655618927473775990157317945366509472028491108236150125473392848896;
            6'd24: xpb[2] = 256'd2650270597167576494374946251114377773749014290599417289895783102670798848;
            6'd25: xpb[2] = 256'd2760698538716225514973902344910810180988556552707726343641440731948748800;
            6'd26: xpb[2] = 256'd2871126480264874535572858438707242588228098814816035397387098361226698752;
            6'd27: xpb[2] = 256'd2981554421813523556171814532503674995467641076924344451132755990504648704;
            6'd28: xpb[2] = 256'd3091982363362172576770770626300107402707183339032653504878413619782598656;
            6'd29: xpb[2] = 256'd3202410304910821597369726720096539809946725601140962558624071249060548608;
            6'd30: xpb[2] = 256'd3312838246459470617968682813892972217186267863249271612369728878338498560;
            6'd31: xpb[2] = 256'd3423266188008119638567638907689404624425810125357580666115386507616448512;
            6'd32: xpb[2] = 256'd3533694129556768659166595001485837031665352387465889719861044136894398464;
            6'd33: xpb[2] = 256'd3644122071105417679765551095282269438904894649574198773606701766172348416;
            6'd34: xpb[2] = 256'd3754550012654066700364507189078701846144436911682507827352359395450298368;
            6'd35: xpb[2] = 256'd3864977954202715720963463282875134253383979173790816881098017024728248320;
            6'd36: xpb[2] = 256'd3975405895751364741562419376671566660623521435899125934843674654006198272;
            6'd37: xpb[2] = 256'd4085833837300013762161375470467999067863063698007434988589332283284148224;
            6'd38: xpb[2] = 256'd4196261778848662782760331564264431475102605960115744042334989912562098176;
            6'd39: xpb[2] = 256'd4306689720397311803359287658060863882342148222224053096080647541840048128;
            6'd40: xpb[2] = 256'd4417117661945960823958243751857296289581690484332362149826305171117998080;
            6'd41: xpb[2] = 256'd4527545603494609844557199845653728696821232746440671203571962800395948032;
            6'd42: xpb[2] = 256'd4637973545043258865156155939450161104060775008548980257317620429673897984;
            6'd43: xpb[2] = 256'd4748401486591907885755112033246593511300317270657289311063278058951847936;
            6'd44: xpb[2] = 256'd4858829428140556906354068127043025918539859532765598364808935688229797888;
            6'd45: xpb[2] = 256'd4969257369689205926953024220839458325779401794873907418554593317507747840;
            6'd46: xpb[2] = 256'd5079685311237854947551980314635890733018944056982216472300250946785697792;
            6'd47: xpb[2] = 256'd5190113252786503968150936408432323140258486319090525526045908576063647744;
            6'd48: xpb[2] = 256'd5300541194335152988749892502228755547498028581198834579791566205341597696;
            6'd49: xpb[2] = 256'd5410969135883802009348848596025187954737570843307143633537223834619547648;
            6'd50: xpb[2] = 256'd5521397077432451029947804689821620361977113105415452687282881463897497600;
            6'd51: xpb[2] = 256'd5631825018981100050546760783618052769216655367523761741028539093175447552;
            6'd52: xpb[2] = 256'd5742252960529749071145716877414485176456197629632070794774196722453397504;
            6'd53: xpb[2] = 256'd5852680902078398091744672971210917583695739891740379848519854351731347456;
            6'd54: xpb[2] = 256'd5963108843627047112343629065007349990935282153848688902265511981009297408;
            6'd55: xpb[2] = 256'd6073536785175696132942585158803782398174824415956997956011169610287247360;
            6'd56: xpb[2] = 256'd6183964726724345153541541252600214805414366678065307009756827239565197312;
            6'd57: xpb[2] = 256'd6294392668272994174140497346396647212653908940173616063502484868843147264;
            6'd58: xpb[2] = 256'd6404820609821643194739453440193079619893451202281925117248142498121097216;
            6'd59: xpb[2] = 256'd6515248551370292215338409533989512027132993464390234170993800127399047168;
            6'd60: xpb[2] = 256'd6625676492918941235937365627785944434372535726498543224739457756676997120;
            6'd61: xpb[2] = 256'd6736104434467590256536321721582376841612077988606852278485115385954947072;
            6'd62: xpb[2] = 256'd6846532376016239277135277815378809248851620250715161332230773015232897024;
            6'd63: xpb[2] = 256'd6956960317564888297734233909175241656091162512823470385976430644510846976;
        endcase
    end

    always_comb begin
        case(flag[3])
            6'd0: xpb[3] = 256'd0;
            6'd1: xpb[3] = 256'd1766847064778384329583297500742918515832676193732944859930522068447199232;
            6'd2: xpb[3] = 256'd3533694129556768659166595001485837031665352387465889719861044136894398464;
            6'd3: xpb[3] = 256'd5300541194335152988749892502228755547498028581198834579791566205341597696;
            6'd4: xpb[3] = 256'd7067388259113537318333190002971674063330704774931779439722088273788796928;
            6'd5: xpb[3] = 256'd8834235323891921647916487503714592579163380968664724299652610342235996160;
            6'd6: xpb[3] = 256'd10601082388670305977499785004457511094996057162397669159583132410683195392;
            6'd7: xpb[3] = 256'd12367929453448690307083082505200429610828733356130614019513654479130394624;
            6'd8: xpb[3] = 256'd14134776518227074636666380005943348126661409549863558879444176547577593856;
            6'd9: xpb[3] = 256'd15901623583005458966249677506686266642494085743596503739374698616024793088;
            6'd10: xpb[3] = 256'd17668470647783843295832975007429185158326761937329448599305220684471992320;
            6'd11: xpb[3] = 256'd19435317712562227625416272508172103674159438131062393459235742752919191552;
            6'd12: xpb[3] = 256'd21202164777340611954999570008915022189992114324795338319166264821366390784;
            6'd13: xpb[3] = 256'd22969011842118996284582867509657940705824790518528283179096786889813590016;
            6'd14: xpb[3] = 256'd24735858906897380614166165010400859221657466712261228039027308958260789248;
            6'd15: xpb[3] = 256'd26502705971675764943749462511143777737490142905994172898957831026707988480;
            6'd16: xpb[3] = 256'd28269553036454149273332760011886696253322819099727117758888353095155187712;
            6'd17: xpb[3] = 256'd30036400101232533602916057512629614769155495293460062618818875163602386944;
            6'd18: xpb[3] = 256'd31803247166010917932499355013372533284988171487193007478749397232049586176;
            6'd19: xpb[3] = 256'd33570094230789302262082652514115451800820847680925952338679919300496785408;
            6'd20: xpb[3] = 256'd35336941295567686591665950014858370316653523874658897198610441368943984640;
            6'd21: xpb[3] = 256'd37103788360346070921249247515601288832486200068391842058540963437391183872;
            6'd22: xpb[3] = 256'd38870635425124455250832545016344207348318876262124786918471485505838383104;
            6'd23: xpb[3] = 256'd40637482489902839580415842517087125864151552455857731778402007574285582336;
            6'd24: xpb[3] = 256'd42404329554681223909999140017830044379984228649590676638332529642732781568;
            6'd25: xpb[3] = 256'd44171176619459608239582437518572962895816904843323621498263051711179980800;
            6'd26: xpb[3] = 256'd45938023684237992569165735019315881411649581037056566358193573779627180032;
            6'd27: xpb[3] = 256'd47704870749016376898749032520058799927482257230789511218124095848074379264;
            6'd28: xpb[3] = 256'd49471717813794761228332330020801718443314933424522456078054617916521578496;
            6'd29: xpb[3] = 256'd51238564878573145557915627521544636959147609618255400937985139984968777728;
            6'd30: xpb[3] = 256'd53005411943351529887498925022287555474980285811988345797915662053415976960;
            6'd31: xpb[3] = 256'd54772259008129914217082222523030473990812962005721290657846184121863176192;
            6'd32: xpb[3] = 256'd56539106072908298546665520023773392506645638199454235517776706190310375424;
            6'd33: xpb[3] = 256'd58305953137686682876248817524516311022478314393187180377707228258757574656;
            6'd34: xpb[3] = 256'd60072800202465067205832115025259229538310990586920125237637750327204773888;
            6'd35: xpb[3] = 256'd61839647267243451535415412526002148054143666780653070097568272395651973120;
            6'd36: xpb[3] = 256'd63606494332021835864998710026745066569976342974386014957498794464099172352;
            6'd37: xpb[3] = 256'd65373341396800220194582007527487985085809019168118959817429316532546371584;
            6'd38: xpb[3] = 256'd67140188461578604524165305028230903601641695361851904677359838600993570816;
            6'd39: xpb[3] = 256'd68907035526356988853748602528973822117474371555584849537290360669440770048;
            6'd40: xpb[3] = 256'd70673882591135373183331900029716740633307047749317794397220882737887969280;
            6'd41: xpb[3] = 256'd72440729655913757512915197530459659149139723943050739257151404806335168512;
            6'd42: xpb[3] = 256'd74207576720692141842498495031202577664972400136783684117081926874782367744;
            6'd43: xpb[3] = 256'd75974423785470526172081792531945496180805076330516628977012448943229566976;
            6'd44: xpb[3] = 256'd77741270850248910501665090032688414696637752524249573836942971011676766208;
            6'd45: xpb[3] = 256'd79508117915027294831248387533431333212470428717982518696873493080123965440;
            6'd46: xpb[3] = 256'd81274964979805679160831685034174251728303104911715463556804015148571164672;
            6'd47: xpb[3] = 256'd83041812044584063490414982534917170244135781105448408416734537217018363904;
            6'd48: xpb[3] = 256'd84808659109362447819998280035660088759968457299181353276665059285465563136;
            6'd49: xpb[3] = 256'd86575506174140832149581577536403007275801133492914298136595581353912762368;
            6'd50: xpb[3] = 256'd88342353238919216479164875037145925791633809686647242996526103422359961600;
            6'd51: xpb[3] = 256'd90109200303697600808748172537888844307466485880380187856456625490807160832;
            6'd52: xpb[3] = 256'd91876047368475985138331470038631762823299162074113132716387147559254360064;
            6'd53: xpb[3] = 256'd93642894433254369467914767539374681339131838267846077576317669627701559296;
            6'd54: xpb[3] = 256'd95409741498032753797498065040117599854964514461579022436248191696148758528;
            6'd55: xpb[3] = 256'd97176588562811138127081362540860518370797190655311967296178713764595957760;
            6'd56: xpb[3] = 256'd98943435627589522456664660041603436886629866849044912156109235833043156992;
            6'd57: xpb[3] = 256'd100710282692367906786247957542346355402462543042777857016039757901490356224;
            6'd58: xpb[3] = 256'd102477129757146291115831255043089273918295219236510801875970279969937555456;
            6'd59: xpb[3] = 256'd104243976821924675445414552543832192434127895430243746735900802038384754688;
            6'd60: xpb[3] = 256'd106010823886703059774997850044575110949960571623976691595831324106831953920;
            6'd61: xpb[3] = 256'd107777670951481444104581147545318029465793247817709636455761846175279153152;
            6'd62: xpb[3] = 256'd109544518016259828434164445046060947981625924011442581315692368243726352384;
            6'd63: xpb[3] = 256'd111311365081038212763747742546803866497458600205175526175622890312173551616;
        endcase
    end

    always_comb begin
        case(flag[4])
            6'd0: xpb[4] = 256'd0;
            6'd1: xpb[4] = 256'd113078212145816597093331040047546785013291276398908471035553412380620750848;
            6'd2: xpb[4] = 256'd226156424291633194186662080095093570026582552797816942071106824761241501696;
            6'd3: xpb[4] = 256'd339234636437449791279993120142640355039873829196725413106660237141862252544;
            6'd4: xpb[4] = 256'd452312848583266388373324160190187140053165105595633884142213649522483003392;
            6'd5: xpb[4] = 256'd565391060729082985466655200237733925066456381994542355177767061903103754240;
            6'd6: xpb[4] = 256'd678469272874899582559986240285280710079747658393450826213320474283724505088;
            6'd7: xpb[4] = 256'd791547485020716179653317280332827495093038934792359297248873886664345255936;
            6'd8: xpb[4] = 256'd904625697166532776746648320380374280106330211191267768284427299044966006784;
            6'd9: xpb[4] = 256'd1017703909312349373839979360427921065119621487590176239319980711425586757632;
            6'd10: xpb[4] = 256'd1130782121458165970933310400475467850132912763989084710355534123806207508480;
            6'd11: xpb[4] = 256'd1243860333603982568026641440523014635146204040387993181391087536186828259328;
            6'd12: xpb[4] = 256'd1356938545749799165119972480570561420159495316786901652426640948567449010176;
            6'd13: xpb[4] = 256'd1470016757895615762213303520618108205172786593185810123462194360948069761024;
            6'd14: xpb[4] = 256'd1583094970041432359306634560665654990186077869584718594497747773328690511872;
            6'd15: xpb[4] = 256'd1696173182187248956399965600713201775199369145983627065533301185709311262720;
            6'd16: xpb[4] = 256'd1809251394333065553493296640760748560212660422382535536568854598089932013568;
            6'd17: xpb[4] = 256'd1922329606478882150586627680808295345225951698781444007604408010470552764416;
            6'd18: xpb[4] = 256'd2035407818624698747679958720855842130239242975180352478639961422851173515264;
            6'd19: xpb[4] = 256'd2148486030770515344773289760903388915252534251579260949675514835231794266112;
            6'd20: xpb[4] = 256'd2261564242916331941866620800950935700265825527978169420711068247612415016960;
            6'd21: xpb[4] = 256'd2374642455062148538959951840998482485279116804377077891746621659993035767808;
            6'd22: xpb[4] = 256'd2487720667207965136053282881046029270292408080775986362782175072373656518656;
            6'd23: xpb[4] = 256'd2600798879353781733146613921093576055305699357174894833817728484754277269504;
            6'd24: xpb[4] = 256'd2713877091499598330239944961141122840318990633573803304853281897134898020352;
            6'd25: xpb[4] = 256'd2826955303645414927333276001188669625332281909972711775888835309515518771200;
            6'd26: xpb[4] = 256'd2940033515791231524426607041236216410345573186371620246924388721896139522048;
            6'd27: xpb[4] = 256'd3053111727937048121519938081283763195358864462770528717959942134276760272896;
            6'd28: xpb[4] = 256'd3166189940082864718613269121331309980372155739169437188995495546657381023744;
            6'd29: xpb[4] = 256'd3279268152228681315706600161378856765385447015568345660031048959038001774592;
            6'd30: xpb[4] = 256'd3392346364374497912799931201426403550398738291967254131066602371418622525440;
            6'd31: xpb[4] = 256'd3505424576520314509893262241473950335412029568366162602102155783799243276288;
            6'd32: xpb[4] = 256'd3618502788666131106986593281521497120425320844765071073137709196179864027136;
            6'd33: xpb[4] = 256'd3731581000811947704079924321569043905438612121163979544173262608560484777984;
            6'd34: xpb[4] = 256'd3844659212957764301173255361616590690451903397562888015208816020941105528832;
            6'd35: xpb[4] = 256'd3957737425103580898266586401664137475465194673961796486244369433321726279680;
            6'd36: xpb[4] = 256'd4070815637249397495359917441711684260478485950360704957279922845702347030528;
            6'd37: xpb[4] = 256'd4183893849395214092453248481759231045491777226759613428315476258082967781376;
            6'd38: xpb[4] = 256'd4296972061541030689546579521806777830505068503158521899351029670463588532224;
            6'd39: xpb[4] = 256'd4410050273686847286639910561854324615518359779557430370386583082844209283072;
            6'd40: xpb[4] = 256'd4523128485832663883733241601901871400531651055956338841422136495224830033920;
            6'd41: xpb[4] = 256'd4636206697978480480826572641949418185544942332355247312457689907605450784768;
            6'd42: xpb[4] = 256'd4749284910124297077919903681996964970558233608754155783493243319986071535616;
            6'd43: xpb[4] = 256'd4862363122270113675013234722044511755571524885153064254528796732366692286464;
            6'd44: xpb[4] = 256'd4975441334415930272106565762092058540584816161551972725564350144747313037312;
            6'd45: xpb[4] = 256'd5088519546561746869199896802139605325598107437950881196599903557127933788160;
            6'd46: xpb[4] = 256'd5201597758707563466293227842187152110611398714349789667635456969508554539008;
            6'd47: xpb[4] = 256'd5314675970853380063386558882234698895624689990748698138671010381889175289856;
            6'd48: xpb[4] = 256'd5427754182999196660479889922282245680637981267147606609706563794269796040704;
            6'd49: xpb[4] = 256'd5540832395145013257573220962329792465651272543546515080742117206650416791552;
            6'd50: xpb[4] = 256'd5653910607290829854666552002377339250664563819945423551777670619031037542400;
            6'd51: xpb[4] = 256'd5766988819436646451759883042424886035677855096344332022813224031411658293248;
            6'd52: xpb[4] = 256'd5880067031582463048853214082472432820691146372743240493848777443792279044096;
            6'd53: xpb[4] = 256'd5993145243728279645946545122519979605704437649142148964884330856172899794944;
            6'd54: xpb[4] = 256'd6106223455874096243039876162567526390717728925541057435919884268553520545792;
            6'd55: xpb[4] = 256'd6219301668019912840133207202615073175731020201939965906955437680934141296640;
            6'd56: xpb[4] = 256'd6332379880165729437226538242662619960744311478338874377990991093314762047488;
            6'd57: xpb[4] = 256'd6445458092311546034319869282710166745757602754737782849026544505695382798336;
            6'd58: xpb[4] = 256'd6558536304457362631413200322757713530770894031136691320062097918076003549184;
            6'd59: xpb[4] = 256'd6671614516603179228506531362805260315784185307535599791097651330456624300032;
            6'd60: xpb[4] = 256'd6784692728748995825599862402852807100797476583934508262133204742837245050880;
            6'd61: xpb[4] = 256'd6897770940894812422693193442900353885810767860333416733168758155217865801728;
            6'd62: xpb[4] = 256'd7010849153040629019786524482947900670824059136732325204204311567598486552576;
            6'd63: xpb[4] = 256'd7123927365186445616879855522995447455837350413131233675239864979979107303424;
        endcase
    end

    always_comb begin
        case(flag[5])
            6'd0: xpb[5] = 256'd0;
            6'd1: xpb[5] = 256'd7237005577332262213973186563042994240850641689530142146275418392359728054272;
            6'd2: xpb[5] = 256'd14474011154664524427946373126085988481701283379060284292550836784719456108544;
            6'd3: xpb[5] = 256'd21711016731996786641919559689128982722551925068590426438826255177079184162816;
            6'd4: xpb[5] = 256'd28948022309329048855892746252171976963402566758120568585101673569438912217088;
            6'd5: xpb[5] = 256'd36185027886661311069865932815214971204253208447650710731377091961798640271360;
            6'd6: xpb[5] = 256'd43422033463993573283839119378257965445103850137180852877652510354158368325632;
            6'd7: xpb[5] = 256'd50659039041325835497812305941300959685954491826710995023927928746518096379904;
            6'd8: xpb[5] = 256'd57896044618658097711785492504343953926805133516241137170203347138877824434176;
            6'd9: xpb[5] = 256'd65133050195990359925758679067386948167655775205771279316478765531237552488448;
            6'd10: xpb[5] = 256'd72370055773322622139731865630429942408506416895301421462754183923597280542720;
            6'd11: xpb[5] = 256'd79607061350654884353705052193472936649357058584831563609029602315957008596992;
            6'd12: xpb[5] = 256'd86844066927987146567678238756515930890207700274361705755305020708316736651264;
            6'd13: xpb[5] = 256'd94081072505319408781651425319558925131058341963891847901580439100676464705536;
            6'd14: xpb[5] = 256'd101318078082651670995624611882601919371908983653421990047855857493036192759808;
            6'd15: xpb[5] = 256'd108555083659983933209597798445644913612759625342952132194131275885395920814080;
            6'd16: xpb[5] = 256'd26959946667150639794667015087359913040558082885985500344465963876353;
            6'd17: xpb[5] = 256'd7237005604292208881123826357710009328210554730088225032260918736825691930625;
            6'd18: xpb[5] = 256'd14474011181624471095097012920753003569061196419618367178536337129185419984897;
            6'd19: xpb[5] = 256'd21711016758956733309070199483795997809911838109148509324811755521545148039169;
            6'd20: xpb[5] = 256'd28948022336288995523043386046838992050762479798678651471087173913904876093441;
            6'd21: xpb[5] = 256'd36185027913621257737016572609881986291613121488208793617362592306264604147713;
            6'd22: xpb[5] = 256'd43422033490953519950989759172924980532463763177738935763638010698624332201985;
            6'd23: xpb[5] = 256'd50659039068285782164962945735967974773314404867269077909913429090984060256257;
            6'd24: xpb[5] = 256'd57896044645618044378936132299010969014165046556799220056188847483343788310529;
            6'd25: xpb[5] = 256'd65133050222950306592909318862053963255015688246329362202464265875703516364801;
            6'd26: xpb[5] = 256'd72370055800282568806882505425096957495866329935859504348739684268063244419073;
            6'd27: xpb[5] = 256'd79607061377614831020855691988139951736716971625389646495015102660422972473345;
            6'd28: xpb[5] = 256'd86844066954947093234828878551182945977567613314919788641290521052782700527617;
            6'd29: xpb[5] = 256'd94081072532279355448802065114225940218418255004449930787565939445142428581889;
            6'd30: xpb[5] = 256'd101318078109611617662775251677268934459268896693980072933841357837502156636161;
            6'd31: xpb[5] = 256'd108555083686943879876748438240311928700119538383510215080116776229861884690433;
            6'd32: xpb[5] = 256'd53919893334301279589334030174719826081116165771971000688931927752706;
            6'd33: xpb[5] = 256'd7237005631252155548274466152377024415570467770646307918246419081291655806978;
            6'd34: xpb[5] = 256'd14474011208584417762247652715420018656421109460176450064521837473651383861250;
            6'd35: xpb[5] = 256'd21711016785916679976220839278463012897271751149706592210797255866011111915522;
            6'd36: xpb[5] = 256'd28948022363248942190194025841506007138122392839236734357072674258370839969794;
            6'd37: xpb[5] = 256'd36185027940581204404167212404549001378973034528766876503348092650730568024066;
            6'd38: xpb[5] = 256'd43422033517913466618140398967591995619823676218297018649623511043090296078338;
            6'd39: xpb[5] = 256'd50659039095245728832113585530634989860674317907827160795898929435450024132610;
            6'd40: xpb[5] = 256'd57896044672577991046086772093677984101524959597357302942174347827809752186882;
            6'd41: xpb[5] = 256'd65133050249910253260059958656720978342375601286887445088449766220169480241154;
            6'd42: xpb[5] = 256'd72370055827242515474033145219763972583226242976417587234725184612529208295426;
            6'd43: xpb[5] = 256'd79607061404574777688006331782806966824076884665947729381000603004888936349698;
            6'd44: xpb[5] = 256'd86844066981907039901979518345849961064927526355477871527276021397248664403970;
            6'd45: xpb[5] = 256'd94081072559239302115952704908892955305778168045008013673551439789608392458242;
            6'd46: xpb[5] = 256'd101318078136571564329925891471935949546628809734538155819826858181968120512514;
            6'd47: xpb[5] = 256'd108555083713903826543899078034978943787479451424068297966102276574327848566786;
            6'd48: xpb[5] = 256'd80879840001451919384001045262079739121674248657956501033397891629059;
            6'd49: xpb[5] = 256'd7237005658212102215425105947044039502930380811204390804231919425757619683331;
            6'd50: xpb[5] = 256'd14474011235544364429398292510087033743781022500734532950507337818117347737603;
            6'd51: xpb[5] = 256'd21711016812876626643371479073130027984631664190264675096782756210477075791875;
            6'd52: xpb[5] = 256'd28948022390208888857344665636173022225482305879794817243058174602836803846147;
            6'd53: xpb[5] = 256'd36185027967541151071317852199216016466332947569324959389333592995196531900419;
            6'd54: xpb[5] = 256'd43422033544873413285291038762259010707183589258855101535609011387556259954691;
            6'd55: xpb[5] = 256'd50659039122205675499264225325302004948034230948385243681884429779915988008963;
            6'd56: xpb[5] = 256'd57896044699537937713237411888344999188884872637915385828159848172275716063235;
            6'd57: xpb[5] = 256'd65133050276870199927210598451387993429735514327445527974435266564635444117507;
            6'd58: xpb[5] = 256'd72370055854202462141183785014430987670586156016975670120710684956995172171779;
            6'd59: xpb[5] = 256'd79607061431534724355156971577473981911436797706505812266986103349354900226051;
            6'd60: xpb[5] = 256'd86844067008866986569130158140516976152287439396035954413261521741714628280323;
            6'd61: xpb[5] = 256'd94081072586199248783103344703559970393138081085566096559536940134074356334595;
            6'd62: xpb[5] = 256'd101318078163531510997076531266602964633988722775096238705812358526434084388867;
            6'd63: xpb[5] = 256'd108555083740863773211049717829645958874839364464626380852087776918793812443139;
        endcase
    end

    always_comb begin
        case(flag[6])
            6'd0: xpb[6] = 256'd0;
            6'd1: xpb[6] = 256'd26959946667150639794667015087359913040558082885985500344465963876353;
            6'd2: xpb[6] = 256'd53919893334301279589334030174719826081116165771971000688931927752706;
            6'd3: xpb[6] = 256'd80879840001451919384001045262079739121674248657956501033397891629059;
            6'd4: xpb[6] = 256'd107839786668602559178668060349439652162232331543942001377863855505412;
            6'd5: xpb[6] = 256'd134799733335753198973335075436799565202790414429927501722329819381765;
            6'd6: xpb[6] = 256'd161759680002903838768002090524159478243348497315913002066795783258118;
            6'd7: xpb[6] = 256'd188719626670054478562669105611519391283906580201898502411261747134471;
            6'd8: xpb[6] = 256'd215679573337205118357336120698879304324464663087884002755727711010824;
            6'd9: xpb[6] = 256'd242639520004355758152003135786239217365022745973869503100193674887177;
            6'd10: xpb[6] = 256'd269599466671506397946670150873599130405580828859855003444659638763530;
            6'd11: xpb[6] = 256'd296559413338657037741337165960959043446138911745840503789125602639883;
            6'd12: xpb[6] = 256'd323519360005807677536004181048318956486696994631826004133591566516236;
            6'd13: xpb[6] = 256'd350479306672958317330671196135678869527255077517811504478057530392589;
            6'd14: xpb[6] = 256'd377439253340108957125338211223038782567813160403797004822523494268942;
            6'd15: xpb[6] = 256'd404399200007259596920005226310398695608371243289782505166989458145295;
            6'd16: xpb[6] = 256'd431359146674410236714672241397758608648929326175768005511455422021648;
            6'd17: xpb[6] = 256'd458319093341560876509339256485118521689487409061753505855921385898001;
            6'd18: xpb[6] = 256'd485279040008711516304006271572478434730045491947739006200387349774354;
            6'd19: xpb[6] = 256'd512238986675862156098673286659838347770603574833724506544853313650707;
            6'd20: xpb[6] = 256'd539198933343012795893340301747198260811161657719710006889319277527060;
            6'd21: xpb[6] = 256'd566158880010163435688007316834558173851719740605695507233785241403413;
            6'd22: xpb[6] = 256'd593118826677314075482674331921918086892277823491681007578251205279766;
            6'd23: xpb[6] = 256'd620078773344464715277341347009277999932835906377666507922717169156119;
            6'd24: xpb[6] = 256'd647038720011615355072008362096637912973393989263652008267183133032472;
            6'd25: xpb[6] = 256'd673998666678765994866675377183997826013952072149637508611649096908825;
            6'd26: xpb[6] = 256'd700958613345916634661342392271357739054510155035623008956115060785178;
            6'd27: xpb[6] = 256'd727918560013067274456009407358717652095068237921608509300581024661531;
            6'd28: xpb[6] = 256'd754878506680217914250676422446077565135626320807594009645046988537884;
            6'd29: xpb[6] = 256'd781838453347368554045343437533437478176184403693579509989512952414237;
            6'd30: xpb[6] = 256'd808798400014519193840010452620797391216742486579565010333978916290590;
            6'd31: xpb[6] = 256'd835758346681669833634677467708157304257300569465550510678444880166943;
            6'd32: xpb[6] = 256'd862718293348820473429344482795517217297858652351536011022910844043296;
            6'd33: xpb[6] = 256'd889678240015971113224011497882877130338416735237521511367376807919649;
            6'd34: xpb[6] = 256'd916638186683121753018678512970237043378974818123507011711842771796002;
            6'd35: xpb[6] = 256'd943598133350272392813345528057596956419532901009492512056308735672355;
            6'd36: xpb[6] = 256'd970558080017423032608012543144956869460090983895478012400774699548708;
            6'd37: xpb[6] = 256'd997518026684573672402679558232316782500649066781463512745240663425061;
            6'd38: xpb[6] = 256'd1024477973351724312197346573319676695541207149667449013089706627301414;
            6'd39: xpb[6] = 256'd1051437920018874951992013588407036608581765232553434513434172591177767;
            6'd40: xpb[6] = 256'd1078397866686025591786680603494396521622323315439420013778638555054120;
            6'd41: xpb[6] = 256'd1105357813353176231581347618581756434662881398325405514123104518930473;
            6'd42: xpb[6] = 256'd1132317760020326871376014633669116347703439481211391014467570482806826;
            6'd43: xpb[6] = 256'd1159277706687477511170681648756476260743997564097376514812036446683179;
            6'd44: xpb[6] = 256'd1186237653354628150965348663843836173784555646983362015156502410559532;
            6'd45: xpb[6] = 256'd1213197600021778790760015678931196086825113729869347515500968374435885;
            6'd46: xpb[6] = 256'd1240157546688929430554682694018555999865671812755333015845434338312238;
            6'd47: xpb[6] = 256'd1267117493356080070349349709105915912906229895641318516189900302188591;
            6'd48: xpb[6] = 256'd1294077440023230710144016724193275825946787978527304016534366266064944;
            6'd49: xpb[6] = 256'd1321037386690381349938683739280635738987346061413289516878832229941297;
            6'd50: xpb[6] = 256'd1347997333357531989733350754367995652027904144299275017223298193817650;
            6'd51: xpb[6] = 256'd1374957280024682629528017769455355565068462227185260517567764157694003;
            6'd52: xpb[6] = 256'd1401917226691833269322684784542715478109020310071246017912230121570356;
            6'd53: xpb[6] = 256'd1428877173358983909117351799630075391149578392957231518256696085446709;
            6'd54: xpb[6] = 256'd1455837120026134548912018814717435304190136475843217018601162049323062;
            6'd55: xpb[6] = 256'd1482797066693285188706685829804795217230694558729202518945628013199415;
            6'd56: xpb[6] = 256'd1509757013360435828501352844892155130271252641615188019290093977075768;
            6'd57: xpb[6] = 256'd1536716960027586468296019859979515043311810724501173519634559940952121;
            6'd58: xpb[6] = 256'd1563676906694737108090686875066874956352368807387159019979025904828474;
            6'd59: xpb[6] = 256'd1590636853361887747885353890154234869392926890273144520323491868704827;
            6'd60: xpb[6] = 256'd1617596800029038387680020905241594782433484973159130020667957832581180;
            6'd61: xpb[6] = 256'd1644556746696189027474687920328954695474043056045115521012423796457533;
            6'd62: xpb[6] = 256'd1671516693363339667269354935416314608514601138931101021356889760333886;
            6'd63: xpb[6] = 256'd1698476640030490307064021950503674521555159221817086521701355724210239;
        endcase
    end

    always_comb begin
        case(flag[7])
            6'd0: xpb[7] = 256'd0;
            6'd1: xpb[7] = 256'd1725436586697640946858688965591034434595717304703072022045821688086592;
            6'd2: xpb[7] = 256'd3450873173395281893717377931182068869191434609406144044091643376173184;
            6'd3: xpb[7] = 256'd5176309760092922840576066896773103303787151914109216066137465064259776;
            6'd4: xpb[7] = 256'd6901746346790563787434755862364137738382869218812288088183286752346368;
            6'd5: xpb[7] = 256'd8627182933488204734293444827955172172978586523515360110229108440432960;
            6'd6: xpb[7] = 256'd10352619520185845681152133793546206607574303828218432132274930128519552;
            6'd7: xpb[7] = 256'd12078056106883486628010822759137241042170021132921504154320751816606144;
            6'd8: xpb[7] = 256'd13803492693581127574869511724728275476765738437624576176366573504692736;
            6'd9: xpb[7] = 256'd15528929280278768521728200690319309911361455742327648198412395192779328;
            6'd10: xpb[7] = 256'd17254365866976409468586889655910344345957173047030720220458216880865920;
            6'd11: xpb[7] = 256'd18979802453674050415445578621501378780552890351733792242504038568952512;
            6'd12: xpb[7] = 256'd20705239040371691362304267587092413215148607656436864264549860257039104;
            6'd13: xpb[7] = 256'd22430675627069332309162956552683447649744324961139936286595681945125696;
            6'd14: xpb[7] = 256'd24156112213766973256021645518274482084340042265843008308641503633212288;
            6'd15: xpb[7] = 256'd25881548800464614202880334483865516518935759570546080330687325321298880;
            6'd16: xpb[7] = 256'd27606985387162255149739023449456550953531476875249152352733147009385472;
            6'd17: xpb[7] = 256'd29332421973859896096597712415047585388127194179952224374778968697472064;
            6'd18: xpb[7] = 256'd31057858560557537043456401380638619822722911484655296396824790385558656;
            6'd19: xpb[7] = 256'd32783295147255177990315090346229654257318628789358368418870612073645248;
            6'd20: xpb[7] = 256'd34508731733952818937173779311820688691914346094061440440916433761731840;
            6'd21: xpb[7] = 256'd36234168320650459884032468277411723126510063398764512462962255449818432;
            6'd22: xpb[7] = 256'd37959604907348100830891157243002757561105780703467584485008077137905024;
            6'd23: xpb[7] = 256'd39685041494045741777749846208593791995701498008170656507053898825991616;
            6'd24: xpb[7] = 256'd41410478080743382724608535174184826430297215312873728529099720514078208;
            6'd25: xpb[7] = 256'd43135914667441023671467224139775860864892932617576800551145542202164800;
            6'd26: xpb[7] = 256'd44861351254138664618325913105366895299488649922279872573191363890251392;
            6'd27: xpb[7] = 256'd46586787840836305565184602070957929734084367226982944595237185578337984;
            6'd28: xpb[7] = 256'd48312224427533946512043291036548964168680084531686016617283007266424576;
            6'd29: xpb[7] = 256'd50037661014231587458901980002139998603275801836389088639328828954511168;
            6'd30: xpb[7] = 256'd51763097600929228405760668967731033037871519141092160661374650642597760;
            6'd31: xpb[7] = 256'd53488534187626869352619357933322067472467236445795232683420472330684352;
            6'd32: xpb[7] = 256'd55213970774324510299478046898913101907062953750498304705466294018770944;
            6'd33: xpb[7] = 256'd56939407361022151246336735864504136341658671055201376727512115706857536;
            6'd34: xpb[7] = 256'd58664843947719792193195424830095170776254388359904448749557937394944128;
            6'd35: xpb[7] = 256'd60390280534417433140054113795686205210850105664607520771603759083030720;
            6'd36: xpb[7] = 256'd62115717121115074086912802761277239645445822969310592793649580771117312;
            6'd37: xpb[7] = 256'd63841153707812715033771491726868274080041540274013664815695402459203904;
            6'd38: xpb[7] = 256'd65566590294510355980630180692459308514637257578716736837741224147290496;
            6'd39: xpb[7] = 256'd67292026881207996927488869658050342949232974883419808859787045835377088;
            6'd40: xpb[7] = 256'd69017463467905637874347558623641377383828692188122880881832867523463680;
            6'd41: xpb[7] = 256'd70742900054603278821206247589232411818424409492825952903878689211550272;
            6'd42: xpb[7] = 256'd72468336641300919768064936554823446253020126797529024925924510899636864;
            6'd43: xpb[7] = 256'd74193773227998560714923625520414480687615844102232096947970332587723456;
            6'd44: xpb[7] = 256'd75919209814696201661782314486005515122211561406935168970016154275810048;
            6'd45: xpb[7] = 256'd77644646401393842608641003451596549556807278711638240992061975963896640;
            6'd46: xpb[7] = 256'd79370082988091483555499692417187583991402996016341313014107797651983232;
            6'd47: xpb[7] = 256'd81095519574789124502358381382778618425998713321044385036153619340069824;
            6'd48: xpb[7] = 256'd82820956161486765449217070348369652860594430625747457058199441028156416;
            6'd49: xpb[7] = 256'd84546392748184406396075759313960687295190147930450529080245262716243008;
            6'd50: xpb[7] = 256'd86271829334882047342934448279551721729785865235153601102291084404329600;
            6'd51: xpb[7] = 256'd87997265921579688289793137245142756164381582539856673124336906092416192;
            6'd52: xpb[7] = 256'd89722702508277329236651826210733790598977299844559745146382727780502784;
            6'd53: xpb[7] = 256'd91448139094974970183510515176324825033573017149262817168428549468589376;
            6'd54: xpb[7] = 256'd93173575681672611130369204141915859468168734453965889190474371156675968;
            6'd55: xpb[7] = 256'd94899012268370252077227893107506893902764451758668961212520192844762560;
            6'd56: xpb[7] = 256'd96624448855067893024086582073097928337360169063372033234566014532849152;
            6'd57: xpb[7] = 256'd98349885441765533970945271038688962771955886368075105256611836220935744;
            6'd58: xpb[7] = 256'd100075322028463174917803960004279997206551603672778177278657657909022336;
            6'd59: xpb[7] = 256'd101800758615160815864662648969871031641147320977481249300703479597108928;
            6'd60: xpb[7] = 256'd103526195201858456811521337935462066075743038282184321322749301285195520;
            6'd61: xpb[7] = 256'd105251631788556097758380026901053100510338755586887393344795122973282112;
            6'd62: xpb[7] = 256'd106977068375253738705238715866644134944934472891590465366840944661368704;
            6'd63: xpb[7] = 256'd108702504961951379652097404832235169379530190196293537388886766349455296;
        endcase
    end

    always_comb begin
        case(flag[8])
            6'd0: xpb[8] = 256'd0;
            6'd1: xpb[8] = 256'd110427941548649020598956093797826203814125907500996609410932588037541888;
            6'd2: xpb[8] = 256'd220855883097298041197912187595652407628251815001993218821865176075083776;
            6'd3: xpb[8] = 256'd331283824645947061796868281393478611442377722502989828232797764112625664;
            6'd4: xpb[8] = 256'd441711766194596082395824375191304815256503630003986437643730352150167552;
            6'd5: xpb[8] = 256'd552139707743245102994780468989131019070629537504983047054662940187709440;
            6'd6: xpb[8] = 256'd662567649291894123593736562786957222884755445005979656465595528225251328;
            6'd7: xpb[8] = 256'd772995590840543144192692656584783426698881352506976265876528116262793216;
            6'd8: xpb[8] = 256'd883423532389192164791648750382609630513007260007972875287460704300335104;
            6'd9: xpb[8] = 256'd993851473937841185390604844180435834327133167508969484698393292337876992;
            6'd10: xpb[8] = 256'd1104279415486490205989560937978262038141259075009966094109325880375418880;
            6'd11: xpb[8] = 256'd1214707357035139226588517031776088241955384982510962703520258468412960768;
            6'd12: xpb[8] = 256'd1325135298583788247187473125573914445769510890011959312931191056450502656;
            6'd13: xpb[8] = 256'd1435563240132437267786429219371740649583636797512955922342123644488044544;
            6'd14: xpb[8] = 256'd1545991181681086288385385313169566853397762705013952531753056232525586432;
            6'd15: xpb[8] = 256'd1656419123229735308984341406967393057211888612514949141163988820563128320;
            6'd16: xpb[8] = 256'd1766847064778384329583297500765219261026014520015945750574921408600670208;
            6'd17: xpb[8] = 256'd1877275006327033350182253594563045464840140427516942359985853996638212096;
            6'd18: xpb[8] = 256'd1987702947875682370781209688360871668654266335017938969396786584675753984;
            6'd19: xpb[8] = 256'd2098130889424331391380165782158697872468392242518935578807719172713295872;
            6'd20: xpb[8] = 256'd2208558830972980411979121875956524076282518150019932188218651760750837760;
            6'd21: xpb[8] = 256'd2318986772521629432578077969754350280096644057520928797629584348788379648;
            6'd22: xpb[8] = 256'd2429414714070278453177034063552176483910769965021925407040516936825921536;
            6'd23: xpb[8] = 256'd2539842655618927473775990157350002687724895872522922016451449524863463424;
            6'd24: xpb[8] = 256'd2650270597167576494374946251147828891539021780023918625862382112901005312;
            6'd25: xpb[8] = 256'd2760698538716225514973902344945655095353147687524915235273314700938547200;
            6'd26: xpb[8] = 256'd2871126480264874535572858438743481299167273595025911844684247288976089088;
            6'd27: xpb[8] = 256'd2981554421813523556171814532541307502981399502526908454095179877013630976;
            6'd28: xpb[8] = 256'd3091982363362172576770770626339133706795525410027905063506112465051172864;
            6'd29: xpb[8] = 256'd3202410304910821597369726720136959910609651317528901672917045053088714752;
            6'd30: xpb[8] = 256'd3312838246459470617968682813934786114423777225029898282327977641126256640;
            6'd31: xpb[8] = 256'd3423266188008119638567638907732612318237903132530894891738910229163798528;
            6'd32: xpb[8] = 256'd3533694129556768659166595001530438522052029040031891501149842817201340416;
            6'd33: xpb[8] = 256'd3644122071105417679765551095328264725866154947532888110560775405238882304;
            6'd34: xpb[8] = 256'd3754550012654066700364507189126090929680280855033884719971707993276424192;
            6'd35: xpb[8] = 256'd3864977954202715720963463282923917133494406762534881329382640581313966080;
            6'd36: xpb[8] = 256'd3975405895751364741562419376721743337308532670035877938793573169351507968;
            6'd37: xpb[8] = 256'd4085833837300013762161375470519569541122658577536874548204505757389049856;
            6'd38: xpb[8] = 256'd4196261778848662782760331564317395744936784485037871157615438345426591744;
            6'd39: xpb[8] = 256'd4306689720397311803359287658115221948750910392538867767026370933464133632;
            6'd40: xpb[8] = 256'd4417117661945960823958243751913048152565036300039864376437303521501675520;
            6'd41: xpb[8] = 256'd4527545603494609844557199845710874356379162207540860985848236109539217408;
            6'd42: xpb[8] = 256'd4637973545043258865156155939508700560193288115041857595259168697576759296;
            6'd43: xpb[8] = 256'd4748401486591907885755112033306526764007414022542854204670101285614301184;
            6'd44: xpb[8] = 256'd4858829428140556906354068127104352967821539930043850814081033873651843072;
            6'd45: xpb[8] = 256'd4969257369689205926953024220902179171635665837544847423491966461689384960;
            6'd46: xpb[8] = 256'd5079685311237854947551980314700005375449791745045844032902899049726926848;
            6'd47: xpb[8] = 256'd5190113252786503968150936408497831579263917652546840642313831637764468736;
            6'd48: xpb[8] = 256'd5300541194335152988749892502295657783078043560047837251724764225802010624;
            6'd49: xpb[8] = 256'd5410969135883802009348848596093483986892169467548833861135696813839552512;
            6'd50: xpb[8] = 256'd5521397077432451029947804689891310190706295375049830470546629401877094400;
            6'd51: xpb[8] = 256'd5631825018981100050546760783689136394520421282550827079957561989914636288;
            6'd52: xpb[8] = 256'd5742252960529749071145716877486962598334547190051823689368494577952178176;
            6'd53: xpb[8] = 256'd5852680902078398091744672971284788802148673097552820298779427165989720064;
            6'd54: xpb[8] = 256'd5963108843627047112343629065082615005962799005053816908190359754027261952;
            6'd55: xpb[8] = 256'd6073536785175696132942585158880441209776924912554813517601292342064803840;
            6'd56: xpb[8] = 256'd6183964726724345153541541252678267413591050820055810127012224930102345728;
            6'd57: xpb[8] = 256'd6294392668272994174140497346476093617405176727556806736423157518139887616;
            6'd58: xpb[8] = 256'd6404820609821643194739453440273919821219302635057803345834090106177429504;
            6'd59: xpb[8] = 256'd6515248551370292215338409534071746025033428542558799955245022694214971392;
            6'd60: xpb[8] = 256'd6625676492918941235937365627869572228847554450059796564655955282252513280;
            6'd61: xpb[8] = 256'd6736104434467590256536321721667398432661680357560793174066887870290055168;
            6'd62: xpb[8] = 256'd6846532376016239277135277815465224636475806265061789783477820458327597056;
            6'd63: xpb[8] = 256'd6956960317564888297734233909263050840289932172562786392888753046365138944;
        endcase
    end

    always_comb begin
        case(flag[9])
            6'd0: xpb[9] = 256'd0;
            6'd1: xpb[9] = 256'd1766847064778384329583297500765219261026014520015945750574921408600670208;
            6'd2: xpb[9] = 256'd3533694129556768659166595001530438522052029040031891501149842817201340416;
            6'd3: xpb[9] = 256'd5300541194335152988749892502295657783078043560047837251724764225802010624;
            6'd4: xpb[9] = 256'd7067388259113537318333190003060877044104058080063783002299685634402680832;
            6'd5: xpb[9] = 256'd8834235323891921647916487503826096305130072600079728752874607043003351040;
            6'd6: xpb[9] = 256'd10601082388670305977499785004591315566156087120095674503449528451604021248;
            6'd7: xpb[9] = 256'd12367929453448690307083082505356534827182101640111620254024449860204691456;
            6'd8: xpb[9] = 256'd14134776518227074636666380006121754088208116160127566004599371268805361664;
            6'd9: xpb[9] = 256'd15901623583005458966249677506886973349234130680143511755174292677406031872;
            6'd10: xpb[9] = 256'd17668470647783843295832975007652192610260145200159457505749214086006702080;
            6'd11: xpb[9] = 256'd19435317712562227625416272508417411871286159720175403256324135494607372288;
            6'd12: xpb[9] = 256'd21202164777340611954999570009182631132312174240191349006899056903208042496;
            6'd13: xpb[9] = 256'd22969011842118996284582867509947850393338188760207294757473978311808712704;
            6'd14: xpb[9] = 256'd24735858906897380614166165010713069654364203280223240508048899720409382912;
            6'd15: xpb[9] = 256'd26502705971675764943749462511478288915390217800239186258623821129010053120;
            6'd16: xpb[9] = 256'd28269553036454149273332760012243508176416232320255132009198742537610723328;
            6'd17: xpb[9] = 256'd30036400101232533602916057513008727437442246840271077759773663946211393536;
            6'd18: xpb[9] = 256'd31803247166010917932499355013773946698468261360287023510348585354812063744;
            6'd19: xpb[9] = 256'd33570094230789302262082652514539165959494275880302969260923506763412733952;
            6'd20: xpb[9] = 256'd35336941295567686591665950015304385220520290400318915011498428172013404160;
            6'd21: xpb[9] = 256'd37103788360346070921249247516069604481546304920334860762073349580614074368;
            6'd22: xpb[9] = 256'd38870635425124455250832545016834823742572319440350806512648270989214744576;
            6'd23: xpb[9] = 256'd40637482489902839580415842517600043003598333960366752263223192397815414784;
            6'd24: xpb[9] = 256'd42404329554681223909999140018365262264624348480382698013798113806416084992;
            6'd25: xpb[9] = 256'd44171176619459608239582437519130481525650363000398643764373035215016755200;
            6'd26: xpb[9] = 256'd45938023684237992569165735019895700786676377520414589514947956623617425408;
            6'd27: xpb[9] = 256'd47704870749016376898749032520660920047702392040430535265522878032218095616;
            6'd28: xpb[9] = 256'd49471717813794761228332330021426139308728406560446481016097799440818765824;
            6'd29: xpb[9] = 256'd51238564878573145557915627522191358569754421080462426766672720849419436032;
            6'd30: xpb[9] = 256'd53005411943351529887498925022956577830780435600478372517247642258020106240;
            6'd31: xpb[9] = 256'd54772259008129914217082222523721797091806450120494318267822563666620776448;
            6'd32: xpb[9] = 256'd56539106072908298546665520024487016352832464640510264018397485075221446656;
            6'd33: xpb[9] = 256'd58305953137686682876248817525252235613858479160526209768972406483822116864;
            6'd34: xpb[9] = 256'd60072800202465067205832115026017454874884493680542155519547327892422787072;
            6'd35: xpb[9] = 256'd61839647267243451535415412526782674135910508200558101270122249301023457280;
            6'd36: xpb[9] = 256'd63606494332021835864998710027547893396936522720574047020697170709624127488;
            6'd37: xpb[9] = 256'd65373341396800220194582007528313112657962537240589992771272092118224797696;
            6'd38: xpb[9] = 256'd67140188461578604524165305029078331918988551760605938521847013526825467904;
            6'd39: xpb[9] = 256'd68907035526356988853748602529843551180014566280621884272421934935426138112;
            6'd40: xpb[9] = 256'd70673882591135373183331900030608770441040580800637830022996856344026808320;
            6'd41: xpb[9] = 256'd72440729655913757512915197531373989702066595320653775773571777752627478528;
            6'd42: xpb[9] = 256'd74207576720692141842498495032139208963092609840669721524146699161228148736;
            6'd43: xpb[9] = 256'd75974423785470526172081792532904428224118624360685667274721620569828818944;
            6'd44: xpb[9] = 256'd77741270850248910501665090033669647485144638880701613025296541978429489152;
            6'd45: xpb[9] = 256'd79508117915027294831248387534434866746170653400717558775871463387030159360;
            6'd46: xpb[9] = 256'd81274964979805679160831685035200086007196667920733504526446384795630829568;
            6'd47: xpb[9] = 256'd83041812044584063490414982535965305268222682440749450277021306204231499776;
            6'd48: xpb[9] = 256'd84808659109362447819998280036730524529248696960765396027596227612832169984;
            6'd49: xpb[9] = 256'd86575506174140832149581577537495743790274711480781341778171149021432840192;
            6'd50: xpb[9] = 256'd88342353238919216479164875038260963051300726000797287528746070430033510400;
            6'd51: xpb[9] = 256'd90109200303697600808748172539026182312326740520813233279320991838634180608;
            6'd52: xpb[9] = 256'd91876047368475985138331470039791401573352755040829179029895913247234850816;
            6'd53: xpb[9] = 256'd93642894433254369467914767540556620834378769560845124780470834655835521024;
            6'd54: xpb[9] = 256'd95409741498032753797498065041321840095404784080861070531045756064436191232;
            6'd55: xpb[9] = 256'd97176588562811138127081362542087059356430798600877016281620677473036861440;
            6'd56: xpb[9] = 256'd98943435627589522456664660042852278617456813120892962032195598881637531648;
            6'd57: xpb[9] = 256'd100710282692367906786247957543617497878482827640908907782770520290238201856;
            6'd58: xpb[9] = 256'd102477129757146291115831255044382717139508842160924853533345441698838872064;
            6'd59: xpb[9] = 256'd104243976821924675445414552545147936400534856680940799283920363107439542272;
            6'd60: xpb[9] = 256'd106010823886703059774997850045913155661560871200956745034495284516040212480;
            6'd61: xpb[9] = 256'd107777670951481444104581147546678374922586885720972690785070205924640882688;
            6'd62: xpb[9] = 256'd109544518016259828434164445047443594183612900240988636535645127333241552896;
            6'd63: xpb[9] = 256'd111311365081038212763747742548208813444638914761004582286220048741842223104;
        endcase
    end

    always_comb begin
        case(flag[10])
            6'd0: xpb[10] = 256'd0;
            6'd1: xpb[10] = 256'd113078212145816597093331040048974032705664929281020528036794970150442893312;
            6'd2: xpb[10] = 256'd226156424291633194186662080097948065411329858562041056073589940300885786624;
            6'd3: xpb[10] = 256'd339234636437449791279993120146922098116994787843061584110384910451328679936;
            6'd4: xpb[10] = 256'd452312848583266388373324160195896130822659717124082112147179880601771573248;
            6'd5: xpb[10] = 256'd565391060729082985466655200244870163528324646405102640183974850752214466560;
            6'd6: xpb[10] = 256'd678469272874899582559986240293844196233989575686123168220769820902657359872;
            6'd7: xpb[10] = 256'd791547485020716179653317280342818228939654504967143696257564791053100253184;
            6'd8: xpb[10] = 256'd904625697166532776746648320391792261645319434248164224294359761203543146496;
            6'd9: xpb[10] = 256'd1017703909312349373839979360440766294350984363529184752331154731353986039808;
            6'd10: xpb[10] = 256'd1130782121458165970933310400489740327056649292810205280367949701504428933120;
            6'd11: xpb[10] = 256'd1243860333603982568026641440538714359762314222091225808404744671654871826432;
            6'd12: xpb[10] = 256'd1356938545749799165119972480587688392467979151372246336441539641805314719744;
            6'd13: xpb[10] = 256'd1470016757895615762213303520636662425173644080653266864478334611955757613056;
            6'd14: xpb[10] = 256'd1583094970041432359306634560685636457879309009934287392515129582106200506368;
            6'd15: xpb[10] = 256'd1696173182187248956399965600734610490584973939215307920551924552256643399680;
            6'd16: xpb[10] = 256'd1809251394333065553493296640783584523290638868496328448588719522407086292992;
            6'd17: xpb[10] = 256'd1922329606478882150586627680832558555996303797777348976625514492557529186304;
            6'd18: xpb[10] = 256'd2035407818624698747679958720881532588701968727058369504662309462707972079616;
            6'd19: xpb[10] = 256'd2148486030770515344773289760930506621407633656339390032699104432858414972928;
            6'd20: xpb[10] = 256'd2261564242916331941866620800979480654113298585620410560735899403008857866240;
            6'd21: xpb[10] = 256'd2374642455062148538959951841028454686818963514901431088772694373159300759552;
            6'd22: xpb[10] = 256'd2487720667207965136053282881077428719524628444182451616809489343309743652864;
            6'd23: xpb[10] = 256'd2600798879353781733146613921126402752230293373463472144846284313460186546176;
            6'd24: xpb[10] = 256'd2713877091499598330239944961175376784935958302744492672883079283610629439488;
            6'd25: xpb[10] = 256'd2826955303645414927333276001224350817641623232025513200919874253761072332800;
            6'd26: xpb[10] = 256'd2940033515791231524426607041273324850347288161306533728956669223911515226112;
            6'd27: xpb[10] = 256'd3053111727937048121519938081322298883052953090587554256993464194061958119424;
            6'd28: xpb[10] = 256'd3166189940082864718613269121371272915758618019868574785030259164212401012736;
            6'd29: xpb[10] = 256'd3279268152228681315706600161420246948464282949149595313067054134362843906048;
            6'd30: xpb[10] = 256'd3392346364374497912799931201469220981169947878430615841103849104513286799360;
            6'd31: xpb[10] = 256'd3505424576520314509893262241518195013875612807711636369140644074663729692672;
            6'd32: xpb[10] = 256'd3618502788666131106986593281567169046581277736992656897177439044814172585984;
            6'd33: xpb[10] = 256'd3731581000811947704079924321616143079286942666273677425214234014964615479296;
            6'd34: xpb[10] = 256'd3844659212957764301173255361665117111992607595554697953251028985115058372608;
            6'd35: xpb[10] = 256'd3957737425103580898266586401714091144698272524835718481287823955265501265920;
            6'd36: xpb[10] = 256'd4070815637249397495359917441763065177403937454116739009324618925415944159232;
            6'd37: xpb[10] = 256'd4183893849395214092453248481812039210109602383397759537361413895566387052544;
            6'd38: xpb[10] = 256'd4296972061541030689546579521861013242815267312678780065398208865716829945856;
            6'd39: xpb[10] = 256'd4410050273686847286639910561909987275520932241959800593435003835867272839168;
            6'd40: xpb[10] = 256'd4523128485832663883733241601958961308226597171240821121471798806017715732480;
            6'd41: xpb[10] = 256'd4636206697978480480826572642007935340932262100521841649508593776168158625792;
            6'd42: xpb[10] = 256'd4749284910124297077919903682056909373637927029802862177545388746318601519104;
            6'd43: xpb[10] = 256'd4862363122270113675013234722105883406343591959083882705582183716469044412416;
            6'd44: xpb[10] = 256'd4975441334415930272106565762154857439049256888364903233618978686619487305728;
            6'd45: xpb[10] = 256'd5088519546561746869199896802203831471754921817645923761655773656769930199040;
            6'd46: xpb[10] = 256'd5201597758707563466293227842252805504460586746926944289692568626920373092352;
            6'd47: xpb[10] = 256'd5314675970853380063386558882301779537166251676207964817729363597070815985664;
            6'd48: xpb[10] = 256'd5427754182999196660479889922350753569871916605488985345766158567221258878976;
            6'd49: xpb[10] = 256'd5540832395145013257573220962399727602577581534770005873802953537371701772288;
            6'd50: xpb[10] = 256'd5653910607290829854666552002448701635283246464051026401839748507522144665600;
            6'd51: xpb[10] = 256'd5766988819436646451759883042497675667988911393332046929876543477672587558912;
            6'd52: xpb[10] = 256'd5880067031582463048853214082546649700694576322613067457913338447823030452224;
            6'd53: xpb[10] = 256'd5993145243728279645946545122595623733400241251894087985950133417973473345536;
            6'd54: xpb[10] = 256'd6106223455874096243039876162644597766105906181175108513986928388123916238848;
            6'd55: xpb[10] = 256'd6219301668019912840133207202693571798811571110456129042023723358274359132160;
            6'd56: xpb[10] = 256'd6332379880165729437226538242742545831517236039737149570060518328424802025472;
            6'd57: xpb[10] = 256'd6445458092311546034319869282791519864222900969018170098097313298575244918784;
            6'd58: xpb[10] = 256'd6558536304457362631413200322840493896928565898299190626134108268725687812096;
            6'd59: xpb[10] = 256'd6671614516603179228506531362889467929634230827580211154170903238876130705408;
            6'd60: xpb[10] = 256'd6784692728748995825599862402938441962339895756861231682207698209026573598720;
            6'd61: xpb[10] = 256'd6897770940894812422693193442987415995045560686142252210244493179177016492032;
            6'd62: xpb[10] = 256'd7010849153040629019786524483036390027751225615423272738281288149327459385344;
            6'd63: xpb[10] = 256'd7123927365186445616879855523085364060456890544704293266318083119477902278656;
        endcase
    end

    always_comb begin
        case(flag[11])
            6'd0: xpb[11] = 256'd0;
            6'd1: xpb[11] = 256'd7237005577332262213973186563134338093162555473985313794354878089628345171968;
            6'd2: xpb[11] = 256'd14474011154664524427946373126268676186325110947970627588709756179256690343936;
            6'd3: xpb[11] = 256'd21711016731996786641919559689403014279487666421955941383064634268885035515904;
            6'd4: xpb[11] = 256'd28948022309329048855892746252537352372650221895941255177419512358513380687872;
            6'd5: xpb[11] = 256'd36185027886661311069865932815671690465812777369926568971774390448141725859840;
            6'd6: xpb[11] = 256'd43422033463993573283839119378806028558975332843911882766129268537770071031808;
            6'd7: xpb[11] = 256'd50659039041325835497812305941940366652137888317897196560484146627398416203776;
            6'd8: xpb[11] = 256'd57896044618658097711785492505074704745300443791882510354839024717026761375744;
            6'd9: xpb[11] = 256'd65133050195990359925758679068209042838462999265867824149193902806655106547712;
            6'd10: xpb[11] = 256'd72370055773322622139731865631343380931625554739853137943548780896283451719680;
            6'd11: xpb[11] = 256'd79607061350654884353705052194477719024788110213838451737903658985911796891648;
            6'd12: xpb[11] = 256'd86844066927987146567678238757612057117950665687823765532258537075540142063616;
            6'd13: xpb[11] = 256'd94081072505319408781651425320746395211113221161809079326613415165168487235584;
            6'd14: xpb[11] = 256'd101318078082651670995624611883880733304275776635794393120968293254796832407552;
            6'd15: xpb[11] = 256'd108555083659983933209597798447015071397438332109779706915323171344425177579520;
            6'd16: xpb[11] = 256'd26959946667150639796128516724350533591840829255256855500763837759489;
            6'd17: xpb[11] = 256'd7237005604292208881123826359262854817513089065826143049611733590392182931457;
            6'd18: xpb[11] = 256'd14474011181624471095097012922397192910675644539811456843966611680020528103425;
            6'd19: xpb[11] = 256'd21711016758956733309070199485531531003838200013796770638321489769648873275393;
            6'd20: xpb[11] = 256'd28948022336288995523043386048665869097000755487782084432676367859277218447361;
            6'd21: xpb[11] = 256'd36185027913621257737016572611800207190163310961767398227031245948905563619329;
            6'd22: xpb[11] = 256'd43422033490953519950989759174934545283325866435752712021386124038533908791297;
            6'd23: xpb[11] = 256'd50659039068285782164962945738068883376488421909738025815741002128162253963265;
            6'd24: xpb[11] = 256'd57896044645618044378936132301203221469650977383723339610095880217790599135233;
            6'd25: xpb[11] = 256'd65133050222950306592909318864337559562813532857708653404450758307418944307201;
            6'd26: xpb[11] = 256'd72370055800282568806882505427471897655976088331693967198805636397047289479169;
            6'd27: xpb[11] = 256'd79607061377614831020855691990606235749138643805679280993160514486675634651137;
            6'd28: xpb[11] = 256'd86844066954947093234828878553740573842301199279664594787515392576303979823105;
            6'd29: xpb[11] = 256'd94081072532279355448802065116874911935463754753649908581870270665932324995073;
            6'd30: xpb[11] = 256'd101318078109611617662775251680009250028626310227635222376225148755560670167041;
            6'd31: xpb[11] = 256'd108555083686943879876748438243143588121788865701620536170580026845189015339009;
            6'd32: xpb[11] = 256'd53919893334301279592257033448701067183681658510513711001527675518978;
            6'd33: xpb[11] = 256'd7237005631252155548274466155391371541863622657666972304868589091156020690946;
            6'd34: xpb[11] = 256'd14474011208584417762247652718525709635026178131652286099223467180784365862914;
            6'd35: xpb[11] = 256'd21711016785916679976220839281660047728188733605637599893578345270412711034882;
            6'd36: xpb[11] = 256'd28948022363248942190194025844794385821351289079622913687933223360041056206850;
            6'd37: xpb[11] = 256'd36185027940581204404167212407928723914513844553608227482288101449669401378818;
            6'd38: xpb[11] = 256'd43422033517913466618140398971063062007676400027593541276642979539297746550786;
            6'd39: xpb[11] = 256'd50659039095245728832113585534197400100838955501578855070997857628926091722754;
            6'd40: xpb[11] = 256'd57896044672577991046086772097331738194001510975564168865352735718554436894722;
            6'd41: xpb[11] = 256'd65133050249910253260059958660466076287164066449549482659707613808182782066690;
            6'd42: xpb[11] = 256'd72370055827242515474033145223600414380326621923534796454062491897811127238658;
            6'd43: xpb[11] = 256'd79607061404574777688006331786734752473489177397520110248417369987439472410626;
            6'd44: xpb[11] = 256'd86844066981907039901979518349869090566651732871505424042772248077067817582594;
            6'd45: xpb[11] = 256'd94081072559239302115952704913003428659814288345490737837127126166696162754562;
            6'd46: xpb[11] = 256'd101318078136571564329925891476137766752976843819476051631482004256324507926530;
            6'd47: xpb[11] = 256'd108555083713903826543899078039272104846139399293461365425836882345952853098498;
            6'd48: xpb[11] = 256'd80879840001451919388385550173051600775522487765770566502291513278467;
            6'd49: xpb[11] = 256'd7237005658212102215425105951519888266214156249507801560125444591919858450435;
            6'd50: xpb[11] = 256'd14474011235544364429398292514654226359376711723493115354480322681548203622403;
            6'd51: xpb[11] = 256'd21711016812876626643371479077788564452539267197478429148835200771176548794371;
            6'd52: xpb[11] = 256'd28948022390208888857344665640922902545701822671463742943190078860804893966339;
            6'd53: xpb[11] = 256'd36185027967541151071317852204057240638864378145449056737544956950433239138307;
            6'd54: xpb[11] = 256'd43422033544873413285291038767191578732026933619434370531899835040061584310275;
            6'd55: xpb[11] = 256'd50659039122205675499264225330325916825189489093419684326254713129689929482243;
            6'd56: xpb[11] = 256'd57896044699537937713237411893460254918352044567404998120609591219318274654211;
            6'd57: xpb[11] = 256'd65133050276870199927210598456594593011514600041390311914964469308946619826179;
            6'd58: xpb[11] = 256'd72370055854202462141183785019728931104677155515375625709319347398574964998147;
            6'd59: xpb[11] = 256'd79607061431534724355156971582863269197839710989360939503674225488203310170115;
            6'd60: xpb[11] = 256'd86844067008866986569130158145997607291002266463346253298029103577831655342083;
            6'd61: xpb[11] = 256'd94081072586199248783103344709131945384164821937331567092383981667460000514051;
            6'd62: xpb[11] = 256'd101318078163531510997076531272266283477327377411316880886738859757088345686019;
            6'd63: xpb[11] = 256'd108555083740863773211049717835400621570489932885302194681093737846716690857987;
        endcase
    end

    always_comb begin
        case(flag[12])
            6'd0: xpb[12] = 256'd0;
            6'd1: xpb[12] = 256'd26959946667150639796128516724350533591840829255256855500763837759489;
            6'd2: xpb[12] = 256'd53919893334301279592257033448701067183681658510513711001527675518978;
            6'd3: xpb[12] = 256'd80879840001451919388385550173051600775522487765770566502291513278467;
            6'd4: xpb[12] = 256'd107839786668602559184514066897402134367363317021027422003055351037956;
            6'd5: xpb[12] = 256'd134799733335753198980642583621752667959204146276284277503819188797445;
            6'd6: xpb[12] = 256'd161759680002903838776771100346103201551044975531541133004583026556934;
            6'd7: xpb[12] = 256'd188719626670054478572899617070453735142885804786797988505346864316423;
            6'd8: xpb[12] = 256'd215679573337205118369028133794804268734726634042054844006110702075912;
            6'd9: xpb[12] = 256'd242639520004355758165156650519154802326567463297311699506874539835401;
            6'd10: xpb[12] = 256'd269599466671506397961285167243505335918408292552568555007638377594890;
            6'd11: xpb[12] = 256'd296559413338657037757413683967855869510249121807825410508402215354379;
            6'd12: xpb[12] = 256'd323519360005807677553542200692206403102089951063082266009166053113868;
            6'd13: xpb[12] = 256'd350479306672958317349670717416556936693930780318339121509929890873357;
            6'd14: xpb[12] = 256'd377439253340108957145799234140907470285771609573595977010693728632846;
            6'd15: xpb[12] = 256'd404399200007259596941927750865258003877612438828852832511457566392335;
            6'd16: xpb[12] = 256'd431359146674410236738056267589608537469453268084109688012221404151824;
            6'd17: xpb[12] = 256'd458319093341560876534184784313959071061294097339366543512985241911313;
            6'd18: xpb[12] = 256'd485279040008711516330313301038309604653134926594623399013749079670802;
            6'd19: xpb[12] = 256'd512238986675862156126441817762660138244975755849880254514512917430291;
            6'd20: xpb[12] = 256'd539198933343012795922570334487010671836816585105137110015276755189780;
            6'd21: xpb[12] = 256'd566158880010163435718698851211361205428657414360393965516040592949269;
            6'd22: xpb[12] = 256'd593118826677314075514827367935711739020498243615650821016804430708758;
            6'd23: xpb[12] = 256'd620078773344464715310955884660062272612339072870907676517568268468247;
            6'd24: xpb[12] = 256'd647038720011615355107084401384412806204179902126164532018332106227736;
            6'd25: xpb[12] = 256'd673998666678765994903212918108763339796020731381421387519095943987225;
            6'd26: xpb[12] = 256'd700958613345916634699341434833113873387861560636678243019859781746714;
            6'd27: xpb[12] = 256'd727918560013067274495469951557464406979702389891935098520623619506203;
            6'd28: xpb[12] = 256'd754878506680217914291598468281814940571543219147191954021387457265692;
            6'd29: xpb[12] = 256'd781838453347368554087726985006165474163384048402448809522151295025181;
            6'd30: xpb[12] = 256'd808798400014519193883855501730516007755224877657705665022915132784670;
            6'd31: xpb[12] = 256'd835758346681669833679984018454866541347065706912962520523678970544159;
            6'd32: xpb[12] = 256'd862718293348820473476112535179217074938906536168219376024442808303648;
            6'd33: xpb[12] = 256'd889678240015971113272241051903567608530747365423476231525206646063137;
            6'd34: xpb[12] = 256'd916638186683121753068369568627918142122588194678733087025970483822626;
            6'd35: xpb[12] = 256'd943598133350272392864498085352268675714429023933989942526734321582115;
            6'd36: xpb[12] = 256'd970558080017423032660626602076619209306269853189246798027498159341604;
            6'd37: xpb[12] = 256'd997518026684573672456755118800969742898110682444503653528261997101093;
            6'd38: xpb[12] = 256'd1024477973351724312252883635525320276489951511699760509029025834860582;
            6'd39: xpb[12] = 256'd1051437920018874952049012152249670810081792340955017364529789672620071;
            6'd40: xpb[12] = 256'd1078397866686025591845140668974021343673633170210274220030553510379560;
            6'd41: xpb[12] = 256'd1105357813353176231641269185698371877265473999465531075531317348139049;
            6'd42: xpb[12] = 256'd1132317760020326871437397702422722410857314828720787931032081185898538;
            6'd43: xpb[12] = 256'd1159277706687477511233526219147072944449155657976044786532845023658027;
            6'd44: xpb[12] = 256'd1186237653354628151029654735871423478040996487231301642033608861417516;
            6'd45: xpb[12] = 256'd1213197600021778790825783252595774011632837316486558497534372699177005;
            6'd46: xpb[12] = 256'd1240157546688929430621911769320124545224678145741815353035136536936494;
            6'd47: xpb[12] = 256'd1267117493356080070418040286044475078816518974997072208535900374695983;
            6'd48: xpb[12] = 256'd1294077440023230710214168802768825612408359804252329064036664212455472;
            6'd49: xpb[12] = 256'd1321037386690381350010297319493176146000200633507585919537428050214961;
            6'd50: xpb[12] = 256'd1347997333357531989806425836217526679592041462762842775038191887974450;
            6'd51: xpb[12] = 256'd1374957280024682629602554352941877213183882292018099630538955725733939;
            6'd52: xpb[12] = 256'd1401917226691833269398682869666227746775723121273356486039719563493428;
            6'd53: xpb[12] = 256'd1428877173358983909194811386390578280367563950528613341540483401252917;
            6'd54: xpb[12] = 256'd1455837120026134548990939903114928813959404779783870197041247239012406;
            6'd55: xpb[12] = 256'd1482797066693285188787068419839279347551245609039127052542011076771895;
            6'd56: xpb[12] = 256'd1509757013360435828583196936563629881143086438294383908042774914531384;
            6'd57: xpb[12] = 256'd1536716960027586468379325453287980414734927267549640763543538752290873;
            6'd58: xpb[12] = 256'd1563676906694737108175453970012330948326768096804897619044302590050362;
            6'd59: xpb[12] = 256'd1590636853361887747971582486736681481918608926060154474545066427809851;
            6'd60: xpb[12] = 256'd1617596800029038387767711003461032015510449755315411330045830265569340;
            6'd61: xpb[12] = 256'd1644556746696189027563839520185382549102290584570668185546594103328829;
            6'd62: xpb[12] = 256'd1671516693363339667359968036909733082694131413825925041047357941088318;
            6'd63: xpb[12] = 256'd1698476640030490307156096553634083616285972243081181896548121778847807;
        endcase
    end

    always_comb begin
        case(flag[13])
            6'd0: xpb[13] = 256'd0;
            6'd1: xpb[13] = 256'd1725436586697640946952225070358434149877813072336438752048885616607296;
            6'd2: xpb[13] = 256'd3450873173395281893904450140716868299755626144672877504097771233214592;
            6'd3: xpb[13] = 256'd5176309760092922840856675211075302449633439217009316256146656849821888;
            6'd4: xpb[13] = 256'd6901746346790563787808900281433736599511252289345755008195542466429184;
            6'd5: xpb[13] = 256'd8627182933488204734761125351792170749389065361682193760244428083036480;
            6'd6: xpb[13] = 256'd10352619520185845681713350422150604899266878434018632512293313699643776;
            6'd7: xpb[13] = 256'd12078056106883486628665575492509039049144691506355071264342199316251072;
            6'd8: xpb[13] = 256'd13803492693581127575617800562867473199022504578691510016391084932858368;
            6'd9: xpb[13] = 256'd15528929280278768522570025633225907348900317651027948768439970549465664;
            6'd10: xpb[13] = 256'd17254365866976409469522250703584341498778130723364387520488856166072960;
            6'd11: xpb[13] = 256'd18979802453674050416474475773942775648655943795700826272537741782680256;
            6'd12: xpb[13] = 256'd20705239040371691363426700844301209798533756868037265024586627399287552;
            6'd13: xpb[13] = 256'd22430675627069332310378925914659643948411569940373703776635513015894848;
            6'd14: xpb[13] = 256'd24156112213766973257331150985018078098289383012710142528684398632502144;
            6'd15: xpb[13] = 256'd25881548800464614204283376055376512248167196085046581280733284249109440;
            6'd16: xpb[13] = 256'd27606985387162255151235601125734946398045009157383020032782169865716736;
            6'd17: xpb[13] = 256'd29332421973859896098187826196093380547922822229719458784831055482324032;
            6'd18: xpb[13] = 256'd31057858560557537045140051266451814697800635302055897536879941098931328;
            6'd19: xpb[13] = 256'd32783295147255177992092276336810248847678448374392336288928826715538624;
            6'd20: xpb[13] = 256'd34508731733952818939044501407168682997556261446728775040977712332145920;
            6'd21: xpb[13] = 256'd36234168320650459885996726477527117147434074519065213793026597948753216;
            6'd22: xpb[13] = 256'd37959604907348100832948951547885551297311887591401652545075483565360512;
            6'd23: xpb[13] = 256'd39685041494045741779901176618243985447189700663738091297124369181967808;
            6'd24: xpb[13] = 256'd41410478080743382726853401688602419597067513736074530049173254798575104;
            6'd25: xpb[13] = 256'd43135914667441023673805626758960853746945326808410968801222140415182400;
            6'd26: xpb[13] = 256'd44861351254138664620757851829319287896823139880747407553271026031789696;
            6'd27: xpb[13] = 256'd46586787840836305567710076899677722046700952953083846305319911648396992;
            6'd28: xpb[13] = 256'd48312224427533946514662301970036156196578766025420285057368797265004288;
            6'd29: xpb[13] = 256'd50037661014231587461614527040394590346456579097756723809417682881611584;
            6'd30: xpb[13] = 256'd51763097600929228408566752110753024496334392170093162561466568498218880;
            6'd31: xpb[13] = 256'd53488534187626869355518977181111458646212205242429601313515454114826176;
            6'd32: xpb[13] = 256'd55213970774324510302471202251469892796090018314766040065564339731433472;
            6'd33: xpb[13] = 256'd56939407361022151249423427321828326945967831387102478817613225348040768;
            6'd34: xpb[13] = 256'd58664843947719792196375652392186761095845644459438917569662110964648064;
            6'd35: xpb[13] = 256'd60390280534417433143327877462545195245723457531775356321710996581255360;
            6'd36: xpb[13] = 256'd62115717121115074090280102532903629395601270604111795073759882197862656;
            6'd37: xpb[13] = 256'd63841153707812715037232327603262063545479083676448233825808767814469952;
            6'd38: xpb[13] = 256'd65566590294510355984184552673620497695356896748784672577857653431077248;
            6'd39: xpb[13] = 256'd67292026881207996931136777743978931845234709821121111329906539047684544;
            6'd40: xpb[13] = 256'd69017463467905637878089002814337365995112522893457550081955424664291840;
            6'd41: xpb[13] = 256'd70742900054603278825041227884695800144990335965793988834004310280899136;
            6'd42: xpb[13] = 256'd72468336641300919771993452955054234294868149038130427586053195897506432;
            6'd43: xpb[13] = 256'd74193773227998560718945678025412668444745962110466866338102081514113728;
            6'd44: xpb[13] = 256'd75919209814696201665897903095771102594623775182803305090150967130721024;
            6'd45: xpb[13] = 256'd77644646401393842612850128166129536744501588255139743842199852747328320;
            6'd46: xpb[13] = 256'd79370082988091483559802353236487970894379401327476182594248738363935616;
            6'd47: xpb[13] = 256'd81095519574789124506754578306846405044257214399812621346297623980542912;
            6'd48: xpb[13] = 256'd82820956161486765453706803377204839194135027472149060098346509597150208;
            6'd49: xpb[13] = 256'd84546392748184406400659028447563273344012840544485498850395395213757504;
            6'd50: xpb[13] = 256'd86271829334882047347611253517921707493890653616821937602444280830364800;
            6'd51: xpb[13] = 256'd87997265921579688294563478588280141643768466689158376354493166446972096;
            6'd52: xpb[13] = 256'd89722702508277329241515703658638575793646279761494815106542052063579392;
            6'd53: xpb[13] = 256'd91448139094974970188467928728997009943524092833831253858590937680186688;
            6'd54: xpb[13] = 256'd93173575681672611135420153799355444093401905906167692610639823296793984;
            6'd55: xpb[13] = 256'd94899012268370252082372378869713878243279718978504131362688708913401280;
            6'd56: xpb[13] = 256'd96624448855067893029324603940072312393157532050840570114737594530008576;
            6'd57: xpb[13] = 256'd98349885441765533976276829010430746543035345123177008866786480146615872;
            6'd58: xpb[13] = 256'd100075322028463174923229054080789180692913158195513447618835365763223168;
            6'd59: xpb[13] = 256'd101800758615160815870181279151147614842790971267849886370884251379830464;
            6'd60: xpb[13] = 256'd103526195201858456817133504221506048992668784340186325122933136996437760;
            6'd61: xpb[13] = 256'd105251631788556097764085729291864483142546597412522763874982022613045056;
            6'd62: xpb[13] = 256'd106977068375253738711037954362222917292424410484859202627030908229652352;
            6'd63: xpb[13] = 256'd108702504961951379657990179432581351442302223557195641379079793846259648;
        endcase
    end

    always_comb begin
        case(flag[14])
            6'd0: xpb[14] = 256'd0;
            6'd1: xpb[14] = 256'd110427941548649020604942404502939785592180036629532080131128679462866944;
            6'd2: xpb[14] = 256'd220855883097298041209884809005879571184360073259064160262257358925733888;
            6'd3: xpb[14] = 256'd331283824645947061814827213508819356776540109888596240393386038388600832;
            6'd4: xpb[14] = 256'd441711766194596082419769618011759142368720146518128320524514717851467776;
            6'd5: xpb[14] = 256'd552139707743245103024712022514698927960900183147660400655643397314334720;
            6'd6: xpb[14] = 256'd662567649291894123629654427017638713553080219777192480786772076777201664;
            6'd7: xpb[14] = 256'd772995590840543144234596831520578499145260256406724560917900756240068608;
            6'd8: xpb[14] = 256'd883423532389192164839539236023518284737440293036256641049029435702935552;
            6'd9: xpb[14] = 256'd993851473937841185444481640526458070329620329665788721180158115165802496;
            6'd10: xpb[14] = 256'd1104279415486490206049424045029397855921800366295320801311286794628669440;
            6'd11: xpb[14] = 256'd1214707357035139226654366449532337641513980402924852881442415474091536384;
            6'd12: xpb[14] = 256'd1325135298583788247259308854035277427106160439554384961573544153554403328;
            6'd13: xpb[14] = 256'd1435563240132437267864251258538217212698340476183917041704672833017270272;
            6'd14: xpb[14] = 256'd1545991181681086288469193663041156998290520512813449121835801512480137216;
            6'd15: xpb[14] = 256'd1656419123229735309074136067544096783882700549442981201966930191943004160;
            6'd16: xpb[14] = 256'd1766847064778384329679078472047036569474880586072513282098058871405871104;
            6'd17: xpb[14] = 256'd1877275006327033350284020876549976355067060622702045362229187550868738048;
            6'd18: xpb[14] = 256'd1987702947875682370888963281052916140659240659331577442360316230331604992;
            6'd19: xpb[14] = 256'd2098130889424331391493905685555855926251420695961109522491444909794471936;
            6'd20: xpb[14] = 256'd2208558830972980412098848090058795711843600732590641602622573589257338880;
            6'd21: xpb[14] = 256'd2318986772521629432703790494561735497435780769220173682753702268720205824;
            6'd22: xpb[14] = 256'd2429414714070278453308732899064675283027960805849705762884830948183072768;
            6'd23: xpb[14] = 256'd2539842655618927473913675303567615068620140842479237843015959627645939712;
            6'd24: xpb[14] = 256'd2650270597167576494518617708070554854212320879108769923147088307108806656;
            6'd25: xpb[14] = 256'd2760698538716225515123560112573494639804500915738302003278216986571673600;
            6'd26: xpb[14] = 256'd2871126480264874535728502517076434425396680952367834083409345666034540544;
            6'd27: xpb[14] = 256'd2981554421813523556333444921579374210988860988997366163540474345497407488;
            6'd28: xpb[14] = 256'd3091982363362172576938387326082313996581041025626898243671603024960274432;
            6'd29: xpb[14] = 256'd3202410304910821597543329730585253782173221062256430323802731704423141376;
            6'd30: xpb[14] = 256'd3312838246459470618148272135088193567765401098885962403933860383886008320;
            6'd31: xpb[14] = 256'd3423266188008119638753214539591133353357581135515494484064989063348875264;
            6'd32: xpb[14] = 256'd3533694129556768659358156944094073138949761172145026564196117742811742208;
            6'd33: xpb[14] = 256'd3644122071105417679963099348597012924541941208774558644327246422274609152;
            6'd34: xpb[14] = 256'd3754550012654066700568041753099952710134121245404090724458375101737476096;
            6'd35: xpb[14] = 256'd3864977954202715721172984157602892495726301282033622804589503781200343040;
            6'd36: xpb[14] = 256'd3975405895751364741777926562105832281318481318663154884720632460663209984;
            6'd37: xpb[14] = 256'd4085833837300013762382868966608772066910661355292686964851761140126076928;
            6'd38: xpb[14] = 256'd4196261778848662782987811371111711852502841391922219044982889819588943872;
            6'd39: xpb[14] = 256'd4306689720397311803592753775614651638095021428551751125114018499051810816;
            6'd40: xpb[14] = 256'd4417117661945960824197696180117591423687201465181283205245147178514677760;
            6'd41: xpb[14] = 256'd4527545603494609844802638584620531209279381501810815285376275857977544704;
            6'd42: xpb[14] = 256'd4637973545043258865407580989123470994871561538440347365507404537440411648;
            6'd43: xpb[14] = 256'd4748401486591907886012523393626410780463741575069879445638533216903278592;
            6'd44: xpb[14] = 256'd4858829428140556906617465798129350566055921611699411525769661896366145536;
            6'd45: xpb[14] = 256'd4969257369689205927222408202632290351648101648328943605900790575829012480;
            6'd46: xpb[14] = 256'd5079685311237854947827350607135230137240281684958475686031919255291879424;
            6'd47: xpb[14] = 256'd5190113252786503968432293011638169922832461721588007766163047934754746368;
            6'd48: xpb[14] = 256'd5300541194335152989037235416141109708424641758217539846294176614217613312;
            6'd49: xpb[14] = 256'd5410969135883802009642177820644049494016821794847071926425305293680480256;
            6'd50: xpb[14] = 256'd5521397077432451030247120225146989279609001831476604006556433973143347200;
            6'd51: xpb[14] = 256'd5631825018981100050852062629649929065201181868106136086687562652606214144;
            6'd52: xpb[14] = 256'd5742252960529749071457005034152868850793361904735668166818691332069081088;
            6'd53: xpb[14] = 256'd5852680902078398092061947438655808636385541941365200246949820011531948032;
            6'd54: xpb[14] = 256'd5963108843627047112666889843158748421977721977994732327080948690994814976;
            6'd55: xpb[14] = 256'd6073536785175696133271832247661688207569902014624264407212077370457681920;
            6'd56: xpb[14] = 256'd6183964726724345153876774652164627993162082051253796487343206049920548864;
            6'd57: xpb[14] = 256'd6294392668272994174481717056667567778754262087883328567474334729383415808;
            6'd58: xpb[14] = 256'd6404820609821643195086659461170507564346442124512860647605463408846282752;
            6'd59: xpb[14] = 256'd6515248551370292215691601865673447349938622161142392727736592088309149696;
            6'd60: xpb[14] = 256'd6625676492918941236296544270176387135530802197771924807867720767772016640;
            6'd61: xpb[14] = 256'd6736104434467590256901486674679326921122982234401456887998849447234883584;
            6'd62: xpb[14] = 256'd6846532376016239277506429079182266706715162271030988968129978126697750528;
            6'd63: xpb[14] = 256'd6956960317564888298111371483685206492307342307660521048261106806160617472;
        endcase
    end

    always_comb begin
        case(flag[15])
            6'd0: xpb[15] = 256'd0;
            6'd1: xpb[15] = 256'd1766847064778384329679078472047036569474880586072513282098058871405871104;
            6'd2: xpb[15] = 256'd3533694129556768659358156944094073138949761172145026564196117742811742208;
            6'd3: xpb[15] = 256'd5300541194335152989037235416141109708424641758217539846294176614217613312;
            6'd4: xpb[15] = 256'd7067388259113537318716313888188146277899522344290053128392235485623484416;
            6'd5: xpb[15] = 256'd8834235323891921648395392360235182847374402930362566410490294357029355520;
            6'd6: xpb[15] = 256'd10601082388670305978074470832282219416849283516435079692588353228435226624;
            6'd7: xpb[15] = 256'd12367929453448690307753549304329255986324164102507592974686412099841097728;
            6'd8: xpb[15] = 256'd14134776518227074637432627776376292555799044688580106256784470971246968832;
            6'd9: xpb[15] = 256'd15901623583005458967111706248423329125273925274652619538882529842652839936;
            6'd10: xpb[15] = 256'd17668470647783843296790784720470365694748805860725132820980588714058711040;
            6'd11: xpb[15] = 256'd19435317712562227626469863192517402264223686446797646103078647585464582144;
            6'd12: xpb[15] = 256'd21202164777340611956148941664564438833698567032870159385176706456870453248;
            6'd13: xpb[15] = 256'd22969011842118996285828020136611475403173447618942672667274765328276324352;
            6'd14: xpb[15] = 256'd24735858906897380615507098608658511972648328205015185949372824199682195456;
            6'd15: xpb[15] = 256'd26502705971675764945186177080705548542123208791087699231470883071088066560;
            6'd16: xpb[15] = 256'd28269553036454149274865255552752585111598089377160212513568941942493937664;
            6'd17: xpb[15] = 256'd30036400101232533604544334024799621681072969963232725795667000813899808768;
            6'd18: xpb[15] = 256'd31803247166010917934223412496846658250547850549305239077765059685305679872;
            6'd19: xpb[15] = 256'd33570094230789302263902490968893694820022731135377752359863118556711550976;
            6'd20: xpb[15] = 256'd35336941295567686593581569440940731389497611721450265641961177428117422080;
            6'd21: xpb[15] = 256'd37103788360346070923260647912987767958972492307522778924059236299523293184;
            6'd22: xpb[15] = 256'd38870635425124455252939726385034804528447372893595292206157295170929164288;
            6'd23: xpb[15] = 256'd40637482489902839582618804857081841097922253479667805488255354042335035392;
            6'd24: xpb[15] = 256'd42404329554681223912297883329128877667397134065740318770353412913740906496;
            6'd25: xpb[15] = 256'd44171176619459608241976961801175914236872014651812832052451471785146777600;
            6'd26: xpb[15] = 256'd45938023684237992571656040273222950806346895237885345334549530656552648704;
            6'd27: xpb[15] = 256'd47704870749016376901335118745269987375821775823957858616647589527958519808;
            6'd28: xpb[15] = 256'd49471717813794761231014197217317023945296656410030371898745648399364390912;
            6'd29: xpb[15] = 256'd51238564878573145560693275689364060514771536996102885180843707270770262016;
            6'd30: xpb[15] = 256'd53005411943351529890372354161411097084246417582175398462941766142176133120;
            6'd31: xpb[15] = 256'd54772259008129914220051432633458133653721298168247911745039825013582004224;
            6'd32: xpb[15] = 256'd56539106072908298549730511105505170223196178754320425027137883884987875328;
            6'd33: xpb[15] = 256'd58305953137686682879409589577552206792671059340392938309235942756393746432;
            6'd34: xpb[15] = 256'd60072800202465067209088668049599243362145939926465451591334001627799617536;
            6'd35: xpb[15] = 256'd61839647267243451538767746521646279931620820512537964873432060499205488640;
            6'd36: xpb[15] = 256'd63606494332021835868446824993693316501095701098610478155530119370611359744;
            6'd37: xpb[15] = 256'd65373341396800220198125903465740353070570581684682991437628178242017230848;
            6'd38: xpb[15] = 256'd67140188461578604527804981937787389640045462270755504719726237113423101952;
            6'd39: xpb[15] = 256'd68907035526356988857484060409834426209520342856828018001824295984828973056;
            6'd40: xpb[15] = 256'd70673882591135373187163138881881462778995223442900531283922354856234844160;
            6'd41: xpb[15] = 256'd72440729655913757516842217353928499348470104028973044566020413727640715264;
            6'd42: xpb[15] = 256'd74207576720692141846521295825975535917944984615045557848118472599046586368;
            6'd43: xpb[15] = 256'd75974423785470526176200374298022572487419865201118071130216531470452457472;
            6'd44: xpb[15] = 256'd77741270850248910505879452770069609056894745787190584412314590341858328576;
            6'd45: xpb[15] = 256'd79508117915027294835558531242116645626369626373263097694412649213264199680;
            6'd46: xpb[15] = 256'd81274964979805679165237609714163682195844506959335610976510708084670070784;
            6'd47: xpb[15] = 256'd83041812044584063494916688186210718765319387545408124258608766956075941888;
            6'd48: xpb[15] = 256'd84808659109362447824595766658257755334794268131480637540706825827481812992;
            6'd49: xpb[15] = 256'd86575506174140832154274845130304791904269148717553150822804884698887684096;
            6'd50: xpb[15] = 256'd88342353238919216483953923602351828473744029303625664104902943570293555200;
            6'd51: xpb[15] = 256'd90109200303697600813633002074398865043218909889698177387001002441699426304;
            6'd52: xpb[15] = 256'd91876047368475985143312080546445901612693790475770690669099061313105297408;
            6'd53: xpb[15] = 256'd93642894433254369472991159018492938182168671061843203951197120184511168512;
            6'd54: xpb[15] = 256'd95409741498032753802670237490539974751643551647915717233295179055917039616;
            6'd55: xpb[15] = 256'd97176588562811138132349315962587011321118432233988230515393237927322910720;
            6'd56: xpb[15] = 256'd98943435627589522462028394434634047890593312820060743797491296798728781824;
            6'd57: xpb[15] = 256'd100710282692367906791707472906681084460068193406133257079589355670134652928;
            6'd58: xpb[15] = 256'd102477129757146291121386551378728121029543073992205770361687414541540524032;
            6'd59: xpb[15] = 256'd104243976821924675451065629850775157599017954578278283643785473412946395136;
            6'd60: xpb[15] = 256'd106010823886703059780744708322822194168492835164350796925883532284352266240;
            6'd61: xpb[15] = 256'd107777670951481444110423786794869230737967715750423310207981591155758137344;
            6'd62: xpb[15] = 256'd109544518016259828440102865266916267307442596336495823490079650027164008448;
            6'd63: xpb[15] = 256'd111311365081038212769781943738963303876917476922568336772177708898569879552;
        endcase
    end

    always_comb begin
        case(flag[16])
            6'd0: xpb[16] = 256'd0;
            6'd1: xpb[16] = 256'd113078212145816597099461022211010340446392357508640850054275767769975750656;
            6'd2: xpb[16] = 256'd226156424291633194198922044422020680892784715017281700108551535539951501312;
            6'd3: xpb[16] = 256'd339234636437449791298383066633031021339177072525922550162827303309927251968;
            6'd4: xpb[16] = 256'd452312848583266388397844088844041361785569430034563400217103071079903002624;
            6'd5: xpb[16] = 256'd565391060729082985497305111055051702231961787543204250271378838849878753280;
            6'd6: xpb[16] = 256'd678469272874899582596766133266062042678354145051845100325654606619854503936;
            6'd7: xpb[16] = 256'd791547485020716179696227155477072383124746502560485950379930374389830254592;
            6'd8: xpb[16] = 256'd904625697166532776795688177688082723571138860069126800434206142159806005248;
            6'd9: xpb[16] = 256'd1017703909312349373895149199899093064017531217577767650488481909929781755904;
            6'd10: xpb[16] = 256'd1130782121458165970994610222110103404463923575086408500542757677699757506560;
            6'd11: xpb[16] = 256'd1243860333603982568094071244321113744910315932595049350597033445469733257216;
            6'd12: xpb[16] = 256'd1356938545749799165193532266532124085356708290103690200651309213239709007872;
            6'd13: xpb[16] = 256'd1470016757895615762292993288743134425803100647612331050705584981009684758528;
            6'd14: xpb[16] = 256'd1583094970041432359392454310954144766249493005120971900759860748779660509184;
            6'd15: xpb[16] = 256'd1696173182187248956491915333165155106695885362629612750814136516549636259840;
            6'd16: xpb[16] = 256'd1809251394333065553591376355376165447142277720138253600868412284319612010496;
            6'd17: xpb[16] = 256'd1922329606478882150690837377587175787588670077646894450922688052089587761152;
            6'd18: xpb[16] = 256'd2035407818624698747790298399798186128035062435155535300976963819859563511808;
            6'd19: xpb[16] = 256'd2148486030770515344889759422009196468481454792664176151031239587629539262464;
            6'd20: xpb[16] = 256'd2261564242916331941989220444220206808927847150172817001085515355399515013120;
            6'd21: xpb[16] = 256'd2374642455062148539088681466431217149374239507681457851139791123169490763776;
            6'd22: xpb[16] = 256'd2487720667207965136188142488642227489820631865190098701194066890939466514432;
            6'd23: xpb[16] = 256'd2600798879353781733287603510853237830267024222698739551248342658709442265088;
            6'd24: xpb[16] = 256'd2713877091499598330387064533064248170713416580207380401302618426479418015744;
            6'd25: xpb[16] = 256'd2826955303645414927486525555275258511159808937716021251356894194249393766400;
            6'd26: xpb[16] = 256'd2940033515791231524585986577486268851606201295224662101411169962019369517056;
            6'd27: xpb[16] = 256'd3053111727937048121685447599697279192052593652733302951465445729789345267712;
            6'd28: xpb[16] = 256'd3166189940082864718784908621908289532498986010241943801519721497559321018368;
            6'd29: xpb[16] = 256'd3279268152228681315884369644119299872945378367750584651573997265329296769024;
            6'd30: xpb[16] = 256'd3392346364374497912983830666330310213391770725259225501628273033099272519680;
            6'd31: xpb[16] = 256'd3505424576520314510083291688541320553838163082767866351682548800869248270336;
            6'd32: xpb[16] = 256'd3618502788666131107182752710752330894284555440276507201736824568639224020992;
            6'd33: xpb[16] = 256'd3731581000811947704282213732963341234730947797785148051791100336409199771648;
            6'd34: xpb[16] = 256'd3844659212957764301381674755174351575177340155293788901845376104179175522304;
            6'd35: xpb[16] = 256'd3957737425103580898481135777385361915623732512802429751899651871949151272960;
            6'd36: xpb[16] = 256'd4070815637249397495580596799596372256070124870311070601953927639719127023616;
            6'd37: xpb[16] = 256'd4183893849395214092680057821807382596516517227819711452008203407489102774272;
            6'd38: xpb[16] = 256'd4296972061541030689779518844018392936962909585328352302062479175259078524928;
            6'd39: xpb[16] = 256'd4410050273686847286878979866229403277409301942836993152116754943029054275584;
            6'd40: xpb[16] = 256'd4523128485832663883978440888440413617855694300345634002171030710799030026240;
            6'd41: xpb[16] = 256'd4636206697978480481077901910651423958302086657854274852225306478569005776896;
            6'd42: xpb[16] = 256'd4749284910124297078177362932862434298748479015362915702279582246338981527552;
            6'd43: xpb[16] = 256'd4862363122270113675276823955073444639194871372871556552333858014108957278208;
            6'd44: xpb[16] = 256'd4975441334415930272376284977284454979641263730380197402388133781878933028864;
            6'd45: xpb[16] = 256'd5088519546561746869475745999495465320087656087888838252442409549648908779520;
            6'd46: xpb[16] = 256'd5201597758707563466575207021706475660534048445397479102496685317418884530176;
            6'd47: xpb[16] = 256'd5314675970853380063674668043917486000980440802906119952550961085188860280832;
            6'd48: xpb[16] = 256'd5427754182999196660774129066128496341426833160414760802605236852958836031488;
            6'd49: xpb[16] = 256'd5540832395145013257873590088339506681873225517923401652659512620728811782144;
            6'd50: xpb[16] = 256'd5653910607290829854973051110550517022319617875432042502713788388498787532800;
            6'd51: xpb[16] = 256'd5766988819436646452072512132761527362766010232940683352768064156268763283456;
            6'd52: xpb[16] = 256'd5880067031582463049171973154972537703212402590449324202822339924038739034112;
            6'd53: xpb[16] = 256'd5993145243728279646271434177183548043658794947957965052876615691808714784768;
            6'd54: xpb[16] = 256'd6106223455874096243370895199394558384105187305466605902930891459578690535424;
            6'd55: xpb[16] = 256'd6219301668019912840470356221605568724551579662975246752985167227348666286080;
            6'd56: xpb[16] = 256'd6332379880165729437569817243816579064997972020483887603039442995118642036736;
            6'd57: xpb[16] = 256'd6445458092311546034669278266027589405444364377992528453093718762888617787392;
            6'd58: xpb[16] = 256'd6558536304457362631768739288238599745890756735501169303147994530658593538048;
            6'd59: xpb[16] = 256'd6671614516603179228868200310449610086337149093009810153202270298428569288704;
            6'd60: xpb[16] = 256'd6784692728748995825967661332660620426783541450518451003256546066198545039360;
            6'd61: xpb[16] = 256'd6897770940894812423067122354871630767229933808027091853310821833968520790016;
            6'd62: xpb[16] = 256'd7010849153040629020166583377082641107676326165535732703365097601738496540672;
            6'd63: xpb[16] = 256'd7123927365186445617266044399293651448122718523044373553419373369508472291328;
        endcase
    end

    always_comb begin
        case(flag[17])
            6'd0: xpb[17] = 256'd0;
            6'd1: xpb[17] = 256'd7237005577332262214365505421504661788569110880553014403473649137278448041984;
            6'd2: xpb[17] = 256'd14474011154664524428731010843009323577138221761106028806947298274556896083968;
            6'd3: xpb[17] = 256'd21711016731996786643096516264513985365707332641659043210420947411835344125952;
            6'd4: xpb[17] = 256'd28948022309329048857462021686018647154276443522212057613894596549113792167936;
            6'd5: xpb[17] = 256'd36185027886661311071827527107523308942845554402765072017368245686392240209920;
            6'd6: xpb[17] = 256'd43422033463993573286193032529027970731414665283318086420841894823670688251904;
            6'd7: xpb[17] = 256'd50659039041325835500558537950532632519983776163871100824315543960949136293888;
            6'd8: xpb[17] = 256'd57896044618658097714924043372037294308552887044424115227789193098227584335872;
            6'd9: xpb[17] = 256'd65133050195990359929289548793541956097121997924977129631262842235506032377856;
            6'd10: xpb[17] = 256'd72370055773322622143655054215046617885691108805530144034736491372784480419840;
            6'd11: xpb[17] = 256'd79607061350654884358020559636551279674260219686083158438210140510062928461824;
            6'd12: xpb[17] = 256'd86844066927987146572386065058055941462829330566636172841683789647341376503808;
            6'd13: xpb[17] = 256'd94081072505319408786751570479560603251398441447189187245157438784619824545792;
            6'd14: xpb[17] = 256'd101318078082651671001117075901065265039967552327742201648631087921898272587776;
            6'd15: xpb[17] = 256'd108555083659983933215482581322569926828536663208295216052104737059176720629760;
            6'd16: xpb[17] = 256'd26959946673427741530053695850855420096924039001157192263165483679745;
            6'd17: xpb[17] = 256'd7237005604292208887793246951558357639424530977477053404630841400443931721729;
            6'd18: xpb[17] = 256'd14474011181624471102158752373063019427993641858030067808104490537722379763713;
            6'd19: xpb[17] = 256'd21711016758956733316524257794567681216562752738583082211578139675000827805697;
            6'd20: xpb[17] = 256'd28948022336288995530889763216072343005131863619136096615051788812279275847681;
            6'd21: xpb[17] = 256'd36185027913621257745255268637577004793700974499689111018525437949557723889665;
            6'd22: xpb[17] = 256'd43422033490953519959620774059081666582270085380242125421999087086836171931649;
            6'd23: xpb[17] = 256'd50659039068285782173986279480586328370839196260795139825472736224114619973633;
            6'd24: xpb[17] = 256'd57896044645618044388351784902090990159408307141348154228946385361393068015617;
            6'd25: xpb[17] = 256'd65133050222950306602717290323595651947977418021901168632420034498671516057601;
            6'd26: xpb[17] = 256'd72370055800282568817082795745100313736546528902454183035893683635949964099585;
            6'd27: xpb[17] = 256'd79607061377614831031448301166604975525115639783007197439367332773228412141569;
            6'd28: xpb[17] = 256'd86844066954947093245813806588109637313684750663560211842840981910506860183553;
            6'd29: xpb[17] = 256'd94081072532279355460179312009614299102253861544113226246314631047785308225537;
            6'd30: xpb[17] = 256'd101318078109611617674544817431118960890822972424666240649788280185063756267521;
            6'd31: xpb[17] = 256'd108555083686943879888910322852623622679392083305219255053261929322342204309505;
            6'd32: xpb[17] = 256'd53919893346855483060107391701710840193848078002314384526330967359490;
            6'd33: xpb[17] = 256'd7237005631252155561220988481612053490279951074401092405788033663609415401474;
            6'd34: xpb[17] = 256'd14474011208584417775586493903116715278849061954954106809261682800887863443458;
            6'd35: xpb[17] = 256'd21711016785916679989951999324621377067418172835507121212735331938166311485442;
            6'd36: xpb[17] = 256'd28948022363248942204317504746126038855987283716060135616208981075444759527426;
            6'd37: xpb[17] = 256'd36185027940581204418683010167630700644556394596613150019682630212723207569410;
            6'd38: xpb[17] = 256'd43422033517913466633048515589135362433125505477166164423156279350001655611394;
            6'd39: xpb[17] = 256'd50659039095245728847414021010640024221694616357719178826629928487280103653378;
            6'd40: xpb[17] = 256'd57896044672577991061779526432144686010263727238272193230103577624558551695362;
            6'd41: xpb[17] = 256'd65133050249910253276145031853649347798832838118825207633577226761836999737346;
            6'd42: xpb[17] = 256'd72370055827242515490510537275154009587401948999378222037050875899115447779330;
            6'd43: xpb[17] = 256'd79607061404574777704876042696658671375971059879931236440524525036393895821314;
            6'd44: xpb[17] = 256'd86844066981907039919241548118163333164540170760484250843998174173672343863298;
            6'd45: xpb[17] = 256'd94081072559239302133607053539667994953109281641037265247471823310950791905282;
            6'd46: xpb[17] = 256'd101318078136571564347972558961172656741678392521590279650945472448229239947266;
            6'd47: xpb[17] = 256'd108555083713903826562338064382677318530247503402143294054419121585507687989250;
            6'd48: xpb[17] = 256'd80879840020283224590161087552566260290772117003471576789496451039235;
            6'd49: xpb[17] = 256'd7237005658212102234648730011665749341135371171325131406945225926774899081219;
            6'd50: xpb[17] = 256'd14474011235544364449014235433170411129704482051878145810418875064053347123203;
            6'd51: xpb[17] = 256'd21711016812876626663379740854675072918273592932431160213892524201331795165187;
            6'd52: xpb[17] = 256'd28948022390208888877745246276179734706842703812984174617366173338610243207171;
            6'd53: xpb[17] = 256'd36185027967541151092110751697684396495411814693537189020839822475888691249155;
            6'd54: xpb[17] = 256'd43422033544873413306476257119189058283980925574090203424313471613167139291139;
            6'd55: xpb[17] = 256'd50659039122205675520841762540693720072550036454643217827787120750445587333123;
            6'd56: xpb[17] = 256'd57896044699537937735207267962198381861119147335196232231260769887724035375107;
            6'd57: xpb[17] = 256'd65133050276870199949572773383703043649688258215749246634734419025002483417091;
            6'd58: xpb[17] = 256'd72370055854202462163938278805207705438257369096302261038208068162280931459075;
            6'd59: xpb[17] = 256'd79607061431534724378303784226712367226826479976855275441681717299559379501059;
            6'd60: xpb[17] = 256'd86844067008866986592669289648217029015395590857408289845155366436837827543043;
            6'd61: xpb[17] = 256'd94081072586199248807034795069721690803964701737961304248629015574116275585027;
            6'd62: xpb[17] = 256'd101318078163531511021400300491226352592533812618514318652102664711394723627011;
            6'd63: xpb[17] = 256'd108555083740863773235765805912731014381102923499067333055576313848673171668995;
        endcase
    end

    always_comb begin
        case(flag[18])
            6'd0: xpb[18] = 256'd0;
            6'd1: xpb[18] = 256'd26959946673427741530053695850855420096924039001157192263165483679745;
            6'd2: xpb[18] = 256'd53919893346855483060107391701710840193848078002314384526330967359490;
            6'd3: xpb[18] = 256'd80879840020283224590161087552566260290772117003471576789496451039235;
            6'd4: xpb[18] = 256'd107839786693710966120214783403421680387696156004628769052661934718980;
            6'd5: xpb[18] = 256'd134799733367138707650268479254277100484620195005785961315827418398725;
            6'd6: xpb[18] = 256'd161759680040566449180322175105132520581544234006943153578992902078470;
            6'd7: xpb[18] = 256'd188719626713994190710375870955987940678468273008100345842158385758215;
            6'd8: xpb[18] = 256'd215679573387421932240429566806843360775392312009257538105323869437960;
            6'd9: xpb[18] = 256'd242639520060849673770483262657698780872316351010414730368489353117705;
            6'd10: xpb[18] = 256'd269599466734277415300536958508554200969240390011571922631654836797450;
            6'd11: xpb[18] = 256'd296559413407705156830590654359409621066164429012729114894820320477195;
            6'd12: xpb[18] = 256'd323519360081132898360644350210265041163088468013886307157985804156940;
            6'd13: xpb[18] = 256'd350479306754560639890698046061120461260012507015043499421151287836685;
            6'd14: xpb[18] = 256'd377439253427988381420751741911975881356936546016200691684316771516430;
            6'd15: xpb[18] = 256'd404399200101416122950805437762831301453860585017357883947482255196175;
            6'd16: xpb[18] = 256'd431359146774843864480859133613686721550784624018515076210647738875920;
            6'd17: xpb[18] = 256'd458319093448271606010912829464542141647708663019672268473813222555665;
            6'd18: xpb[18] = 256'd485279040121699347540966525315397561744632702020829460736978706235410;
            6'd19: xpb[18] = 256'd512238986795127089071020221166252981841556741021986653000144189915155;
            6'd20: xpb[18] = 256'd539198933468554830601073917017108401938480780023143845263309673594900;
            6'd21: xpb[18] = 256'd566158880141982572131127612867963822035404819024301037526475157274645;
            6'd22: xpb[18] = 256'd593118826815410313661181308718819242132328858025458229789640640954390;
            6'd23: xpb[18] = 256'd620078773488838055191235004569674662229252897026615422052806124634135;
            6'd24: xpb[18] = 256'd647038720162265796721288700420530082326176936027772614315971608313880;
            6'd25: xpb[18] = 256'd673998666835693538251342396271385502423100975028929806579137091993625;
            6'd26: xpb[18] = 256'd700958613509121279781396092122240922520025014030086998842302575673370;
            6'd27: xpb[18] = 256'd727918560182549021311449787973096342616949053031244191105468059353115;
            6'd28: xpb[18] = 256'd754878506855976762841503483823951762713873092032401383368633543032860;
            6'd29: xpb[18] = 256'd781838453529404504371557179674807182810797131033558575631799026712605;
            6'd30: xpb[18] = 256'd808798400202832245901610875525662602907721170034715767894964510392350;
            6'd31: xpb[18] = 256'd835758346876259987431664571376518023004645209035872960158129994072095;
            6'd32: xpb[18] = 256'd862718293549687728961718267227373443101569248037030152421295477751840;
            6'd33: xpb[18] = 256'd889678240223115470491771963078228863198493287038187344684460961431585;
            6'd34: xpb[18] = 256'd916638186896543212021825658929084283295417326039344536947626445111330;
            6'd35: xpb[18] = 256'd943598133569970953551879354779939703392341365040501729210791928791075;
            6'd36: xpb[18] = 256'd970558080243398695081933050630795123489265404041658921473957412470820;
            6'd37: xpb[18] = 256'd997518026916826436611986746481650543586189443042816113737122896150565;
            6'd38: xpb[18] = 256'd1024477973590254178142040442332505963683113482043973306000288379830310;
            6'd39: xpb[18] = 256'd1051437920263681919672094138183361383780037521045130498263453863510055;
            6'd40: xpb[18] = 256'd1078397866937109661202147834034216803876961560046287690526619347189800;
            6'd41: xpb[18] = 256'd1105357813610537402732201529885072223973885599047444882789784830869545;
            6'd42: xpb[18] = 256'd1132317760283965144262255225735927644070809638048602075052950314549290;
            6'd43: xpb[18] = 256'd1159277706957392885792308921586783064167733677049759267316115798229035;
            6'd44: xpb[18] = 256'd1186237653630820627322362617437638484264657716050916459579281281908780;
            6'd45: xpb[18] = 256'd1213197600304248368852416313288493904361581755052073651842446765588525;
            6'd46: xpb[18] = 256'd1240157546977676110382470009139349324458505794053230844105612249268270;
            6'd47: xpb[18] = 256'd1267117493651103851912523704990204744555429833054388036368777732948015;
            6'd48: xpb[18] = 256'd1294077440324531593442577400841060164652353872055545228631943216627760;
            6'd49: xpb[18] = 256'd1321037386997959334972631096691915584749277911056702420895108700307505;
            6'd50: xpb[18] = 256'd1347997333671387076502684792542771004846201950057859613158274183987250;
            6'd51: xpb[18] = 256'd1374957280344814818032738488393626424943125989059016805421439667666995;
            6'd52: xpb[18] = 256'd1401917227018242559562792184244481845040050028060173997684605151346740;
            6'd53: xpb[18] = 256'd1428877173691670301092845880095337265136974067061331189947770635026485;
            6'd54: xpb[18] = 256'd1455837120365098042622899575946192685233898106062488382210936118706230;
            6'd55: xpb[18] = 256'd1482797067038525784152953271797048105330822145063645574474101602385975;
            6'd56: xpb[18] = 256'd1509757013711953525683006967647903525427746184064802766737267086065720;
            6'd57: xpb[18] = 256'd1536716960385381267213060663498758945524670223065959959000432569745465;
            6'd58: xpb[18] = 256'd1563676907058809008743114359349614365621594262067117151263598053425210;
            6'd59: xpb[18] = 256'd1590636853732236750273168055200469785718518301068274343526763537104955;
            6'd60: xpb[18] = 256'd1617596800405664491803221751051325205815442340069431535789929020784700;
            6'd61: xpb[18] = 256'd1644556747079092233333275446902180625912366379070588728053094504464445;
            6'd62: xpb[18] = 256'd1671516693752519974863329142753036046009290418071745920316259988144190;
            6'd63: xpb[18] = 256'd1698476640425947716393382838603891466106214457072903112579425471823935;
        endcase
    end

    always_comb begin
        case(flag[19])
            6'd0: xpb[19] = 256'd0;
            6'd1: xpb[19] = 256'd1725436587099375457923436534454746886203138496074060304842590955503680;
            6'd2: xpb[19] = 256'd3450873174198750915846873068909493772406276992148120609685181911007360;
            6'd3: xpb[19] = 256'd5176309761298126373770309603364240658609415488222180914527772866511040;
            6'd4: xpb[19] = 256'd6901746348397501831693746137818987544812553984296241219370363822014720;
            6'd5: xpb[19] = 256'd8627182935496877289617182672273734431015692480370301524212954777518400;
            6'd6: xpb[19] = 256'd10352619522596252747540619206728481317218830976444361829055545733022080;
            6'd7: xpb[19] = 256'd12078056109695628205464055741183228203421969472518422133898136688525760;
            6'd8: xpb[19] = 256'd13803492696795003663387492275637975089625107968592482438740727644029440;
            6'd9: xpb[19] = 256'd15528929283894379121310928810092721975828246464666542743583318599533120;
            6'd10: xpb[19] = 256'd17254365870993754579234365344547468862031384960740603048425909555036800;
            6'd11: xpb[19] = 256'd18979802458093130037157801879002215748234523456814663353268500510540480;
            6'd12: xpb[19] = 256'd20705239045192505495081238413456962634437661952888723658111091466044160;
            6'd13: xpb[19] = 256'd22430675632291880953004674947911709520640800448962783962953682421547840;
            6'd14: xpb[19] = 256'd24156112219391256410928111482366456406843938945036844267796273377051520;
            6'd15: xpb[19] = 256'd25881548806490631868851548016821203293047077441110904572638864332555200;
            6'd16: xpb[19] = 256'd27606985393590007326774984551275950179250215937184964877481455288058880;
            6'd17: xpb[19] = 256'd29332421980689382784698421085730697065453354433259025182324046243562560;
            6'd18: xpb[19] = 256'd31057858567788758242621857620185443951656492929333085487166637199066240;
            6'd19: xpb[19] = 256'd32783295154888133700545294154640190837859631425407145792009228154569920;
            6'd20: xpb[19] = 256'd34508731741987509158468730689094937724062769921481206096851819110073600;
            6'd21: xpb[19] = 256'd36234168329086884616392167223549684610265908417555266401694410065577280;
            6'd22: xpb[19] = 256'd37959604916186260074315603758004431496469046913629326706537001021080960;
            6'd23: xpb[19] = 256'd39685041503285635532239040292459178382672185409703387011379591976584640;
            6'd24: xpb[19] = 256'd41410478090385010990162476826913925268875323905777447316222182932088320;
            6'd25: xpb[19] = 256'd43135914677484386448085913361368672155078462401851507621064773887592000;
            6'd26: xpb[19] = 256'd44861351264583761906009349895823419041281600897925567925907364843095680;
            6'd27: xpb[19] = 256'd46586787851683137363932786430278165927484739393999628230749955798599360;
            6'd28: xpb[19] = 256'd48312224438782512821856222964732912813687877890073688535592546754103040;
            6'd29: xpb[19] = 256'd50037661025881888279779659499187659699891016386147748840435137709606720;
            6'd30: xpb[19] = 256'd51763097612981263737703096033642406586094154882221809145277728665110400;
            6'd31: xpb[19] = 256'd53488534200080639195626532568097153472297293378295869450120319620614080;
            6'd32: xpb[19] = 256'd55213970787180014653549969102551900358500431874369929754962910576117760;
            6'd33: xpb[19] = 256'd56939407374279390111473405637006647244703570370443990059805501531621440;
            6'd34: xpb[19] = 256'd58664843961378765569396842171461394130906708866518050364648092487125120;
            6'd35: xpb[19] = 256'd60390280548478141027320278705916141017109847362592110669490683442628800;
            6'd36: xpb[19] = 256'd62115717135577516485243715240370887903312985858666170974333274398132480;
            6'd37: xpb[19] = 256'd63841153722676891943167151774825634789516124354740231279175865353636160;
            6'd38: xpb[19] = 256'd65566590309776267401090588309280381675719262850814291584018456309139840;
            6'd39: xpb[19] = 256'd67292026896875642859014024843735128561922401346888351888861047264643520;
            6'd40: xpb[19] = 256'd69017463483975018316937461378189875448125539842962412193703638220147200;
            6'd41: xpb[19] = 256'd70742900071074393774860897912644622334328678339036472498546229175650880;
            6'd42: xpb[19] = 256'd72468336658173769232784334447099369220531816835110532803388820131154560;
            6'd43: xpb[19] = 256'd74193773245273144690707770981554116106734955331184593108231411086658240;
            6'd44: xpb[19] = 256'd75919209832372520148631207516008862992938093827258653413074002042161920;
            6'd45: xpb[19] = 256'd77644646419471895606554644050463609879141232323332713717916592997665600;
            6'd46: xpb[19] = 256'd79370083006571271064478080584918356765344370819406774022759183953169280;
            6'd47: xpb[19] = 256'd81095519593670646522401517119373103651547509315480834327601774908672960;
            6'd48: xpb[19] = 256'd82820956180770021980324953653827850537750647811554894632444365864176640;
            6'd49: xpb[19] = 256'd84546392767869397438248390188282597423953786307628954937286956819680320;
            6'd50: xpb[19] = 256'd86271829354968772896171826722737344310156924803703015242129547775184000;
            6'd51: xpb[19] = 256'd87997265942068148354095263257192091196360063299777075546972138730687680;
            6'd52: xpb[19] = 256'd89722702529167523812018699791646838082563201795851135851814729686191360;
            6'd53: xpb[19] = 256'd91448139116266899269942136326101584968766340291925196156657320641695040;
            6'd54: xpb[19] = 256'd93173575703366274727865572860556331854969478787999256461499911597198720;
            6'd55: xpb[19] = 256'd94899012290465650185789009395011078741172617284073316766342502552702400;
            6'd56: xpb[19] = 256'd96624448877565025643712445929465825627375755780147377071185093508206080;
            6'd57: xpb[19] = 256'd98349885464664401101635882463920572513578894276221437376027684463709760;
            6'd58: xpb[19] = 256'd100075322051763776559559318998375319399782032772295497680870275419213440;
            6'd59: xpb[19] = 256'd101800758638863152017482755532830066285985171268369557985712866374717120;
            6'd60: xpb[19] = 256'd103526195225962527475406192067284813172188309764443618290555457330220800;
            6'd61: xpb[19] = 256'd105251631813061902933329628601739560058391448260517678595398048285724480;
            6'd62: xpb[19] = 256'd106977068400161278391253065136194306944594586756591738900240639241228160;
            6'd63: xpb[19] = 256'd108702504987260653849176501670649053830797725252665799205083230196731840;
        endcase
    end

    always_comb begin
        case(flag[20])
            6'd0: xpb[20] = 256'd0;
            6'd1: xpb[20] = 256'd110427941574360029307099938205103800717000863748739859509925821152235520;
            6'd2: xpb[20] = 256'd220855883148720058614199876410207601434001727497479719019851642304471040;
            6'd3: xpb[20] = 256'd331283824723080087921299814615311402151002591246219578529777463456706560;
            6'd4: xpb[20] = 256'd441711766297440117228399752820415202868003454994959438039703284608942080;
            6'd5: xpb[20] = 256'd552139707871800146535499691025519003585004318743699297549629105761177600;
            6'd6: xpb[20] = 256'd662567649446160175842599629230622804302005182492439157059554926913413120;
            6'd7: xpb[20] = 256'd772995591020520205149699567435726605019006046241179016569480748065648640;
            6'd8: xpb[20] = 256'd883423532594880234456799505640830405736006909989918876079406569217884160;
            6'd9: xpb[20] = 256'd993851474169240263763899443845934206453007773738658735589332390370119680;
            6'd10: xpb[20] = 256'd1104279415743600293070999382051038007170008637487398595099258211522355200;
            6'd11: xpb[20] = 256'd1214707357317960322378099320256141807887009501236138454609184032674590720;
            6'd12: xpb[20] = 256'd1325135298892320351685199258461245608604010364984878314119109853826826240;
            6'd13: xpb[20] = 256'd1435563240466680380992299196666349409321011228733618173629035674979061760;
            6'd14: xpb[20] = 256'd1545991182041040410299399134871453210038012092482358033138961496131297280;
            6'd15: xpb[20] = 256'd1656419123615400439606499073076557010755012956231097892648887317283532800;
            6'd16: xpb[20] = 256'd1766847065189760468913599011281660811472013819979837752158813138435768320;
            6'd17: xpb[20] = 256'd1877275006764120498220698949486764612189014683728577611668738959588003840;
            6'd18: xpb[20] = 256'd1987702948338480527527798887691868412906015547477317471178664780740239360;
            6'd19: xpb[20] = 256'd2098130889912840556834898825896972213623016411226057330688590601892474880;
            6'd20: xpb[20] = 256'd2208558831487200586141998764102076014340017274974797190198516423044710400;
            6'd21: xpb[20] = 256'd2318986773061560615449098702307179815057018138723537049708442244196945920;
            6'd22: xpb[20] = 256'd2429414714635920644756198640512283615774019002472276909218368065349181440;
            6'd23: xpb[20] = 256'd2539842656210280674063298578717387416491019866221016768728293886501416960;
            6'd24: xpb[20] = 256'd2650270597784640703370398516922491217208020729969756628238219707653652480;
            6'd25: xpb[20] = 256'd2760698539359000732677498455127595017925021593718496487748145528805888000;
            6'd26: xpb[20] = 256'd2871126480933360761984598393332698818642022457467236347258071349958123520;
            6'd27: xpb[20] = 256'd2981554422507720791291698331537802619359023321215976206767997171110359040;
            6'd28: xpb[20] = 256'd3091982364082080820598798269742906420076024184964716066277922992262594560;
            6'd29: xpb[20] = 256'd3202410305656440849905898207948010220793025048713455925787848813414830080;
            6'd30: xpb[20] = 256'd3312838247230800879212998146153114021510025912462195785297774634567065600;
            6'd31: xpb[20] = 256'd3423266188805160908520098084358217822227026776210935644807700455719301120;
            6'd32: xpb[20] = 256'd3533694130379520937827198022563321622944027639959675504317626276871536640;
            6'd33: xpb[20] = 256'd3644122071953880967134297960768425423661028503708415363827552098023772160;
            6'd34: xpb[20] = 256'd3754550013528240996441397898973529224378029367457155223337477919176007680;
            6'd35: xpb[20] = 256'd3864977955102601025748497837178633025095030231205895082847403740328243200;
            6'd36: xpb[20] = 256'd3975405896676961055055597775383736825812031094954634942357329561480478720;
            6'd37: xpb[20] = 256'd4085833838251321084362697713588840626529031958703374801867255382632714240;
            6'd38: xpb[20] = 256'd4196261779825681113669797651793944427246032822452114661377181203784949760;
            6'd39: xpb[20] = 256'd4306689721400041142976897589999048227963033686200854520887107024937185280;
            6'd40: xpb[20] = 256'd4417117662974401172283997528204152028680034549949594380397032846089420800;
            6'd41: xpb[20] = 256'd4527545604548761201591097466409255829397035413698334239906958667241656320;
            6'd42: xpb[20] = 256'd4637973546123121230898197404614359630114036277447074099416884488393891840;
            6'd43: xpb[20] = 256'd4748401487697481260205297342819463430831037141195813958926810309546127360;
            6'd44: xpb[20] = 256'd4858829429271841289512397281024567231548038004944553818436736130698362880;
            6'd45: xpb[20] = 256'd4969257370846201318819497219229671032265038868693293677946661951850598400;
            6'd46: xpb[20] = 256'd5079685312420561348126597157434774832982039732442033537456587773002833920;
            6'd47: xpb[20] = 256'd5190113253994921377433697095639878633699040596190773396966513594155069440;
            6'd48: xpb[20] = 256'd5300541195569281406740797033844982434416041459939513256476439415307304960;
            6'd49: xpb[20] = 256'd5410969137143641436047896972050086235133042323688253115986365236459540480;
            6'd50: xpb[20] = 256'd5521397078718001465354996910255190035850043187436992975496291057611776000;
            6'd51: xpb[20] = 256'd5631825020292361494662096848460293836567044051185732835006216878764011520;
            6'd52: xpb[20] = 256'd5742252961866721523969196786665397637284044914934472694516142699916247040;
            6'd53: xpb[20] = 256'd5852680903441081553276296724870501438001045778683212554026068521068482560;
            6'd54: xpb[20] = 256'd5963108845015441582583396663075605238718046642431952413535994342220718080;
            6'd55: xpb[20] = 256'd6073536786589801611890496601280709039435047506180692273045920163372953600;
            6'd56: xpb[20] = 256'd6183964728164161641197596539485812840152048369929432132555845984525189120;
            6'd57: xpb[20] = 256'd6294392669738521670504696477690916640869049233678171992065771805677424640;
            6'd58: xpb[20] = 256'd6404820611312881699811796415896020441586050097426911851575697626829660160;
            6'd59: xpb[20] = 256'd6515248552887241729118896354101124242303050961175651711085623447981895680;
            6'd60: xpb[20] = 256'd6625676494461601758425996292306228043020051824924391570595549269134131200;
            6'd61: xpb[20] = 256'd6736104436035961787733096230511331843737052688673131430105475090286366720;
            6'd62: xpb[20] = 256'd6846532377610321817040196168716435644454053552421871289615400911438602240;
            6'd63: xpb[20] = 256'd6956960319184681846347296106921539445171054416170611149125326732590837760;
        endcase
    end

    always_comb begin
        case(flag[21])
            6'd0: xpb[21] = 256'd0;
            6'd1: xpb[21] = 256'd1766847065189760468913599011281660811472013819979837752158813138435768320;
            6'd2: xpb[21] = 256'd3533694130379520937827198022563321622944027639959675504317626276871536640;
            6'd3: xpb[21] = 256'd5300541195569281406740797033844982434416041459939513256476439415307304960;
            6'd4: xpb[21] = 256'd7067388260759041875654396045126643245888055279919351008635252553743073280;
            6'd5: xpb[21] = 256'd8834235325948802344567995056408304057360069099899188760794065692178841600;
            6'd6: xpb[21] = 256'd10601082391138562813481594067689964868832082919879026512952878830614609920;
            6'd7: xpb[21] = 256'd12367929456328323282395193078971625680304096739858864265111691969050378240;
            6'd8: xpb[21] = 256'd14134776521518083751308792090253286491776110559838702017270505107486146560;
            6'd9: xpb[21] = 256'd15901623586707844220222391101534947303248124379818539769429318245921914880;
            6'd10: xpb[21] = 256'd17668470651897604689135990112816608114720138199798377521588131384357683200;
            6'd11: xpb[21] = 256'd19435317717087365158049589124098268926192152019778215273746944522793451520;
            6'd12: xpb[21] = 256'd21202164782277125626963188135379929737664165839758053025905757661229219840;
            6'd13: xpb[21] = 256'd22969011847466886095876787146661590549136179659737890778064570799664988160;
            6'd14: xpb[21] = 256'd24735858912656646564790386157943251360608193479717728530223383938100756480;
            6'd15: xpb[21] = 256'd26502705977846407033703985169224912172080207299697566282382197076536524800;
            6'd16: xpb[21] = 256'd28269553043036167502617584180506572983552221119677404034541010214972293120;
            6'd17: xpb[21] = 256'd30036400108225927971531183191788233795024234939657241786699823353408061440;
            6'd18: xpb[21] = 256'd31803247173415688440444782203069894606496248759637079538858636491843829760;
            6'd19: xpb[21] = 256'd33570094238605448909358381214351555417968262579616917291017449630279598080;
            6'd20: xpb[21] = 256'd35336941303795209378271980225633216229440276399596755043176262768715366400;
            6'd21: xpb[21] = 256'd37103788368984969847185579236914877040912290219576592795335075907151134720;
            6'd22: xpb[21] = 256'd38870635434174730316099178248196537852384304039556430547493889045586903040;
            6'd23: xpb[21] = 256'd40637482499364490785012777259478198663856317859536268299652702184022671360;
            6'd24: xpb[21] = 256'd42404329564554251253926376270759859475328331679516106051811515322458439680;
            6'd25: xpb[21] = 256'd44171176629744011722839975282041520286800345499495943803970328460894208000;
            6'd26: xpb[21] = 256'd45938023694933772191753574293323181098272359319475781556129141599329976320;
            6'd27: xpb[21] = 256'd47704870760123532660667173304604841909744373139455619308287954737765744640;
            6'd28: xpb[21] = 256'd49471717825313293129580772315886502721216386959435457060446767876201512960;
            6'd29: xpb[21] = 256'd51238564890503053598494371327168163532688400779415294812605581014637281280;
            6'd30: xpb[21] = 256'd53005411955692814067407970338449824344160414599395132564764394153073049600;
            6'd31: xpb[21] = 256'd54772259020882574536321569349731485155632428419374970316923207291508817920;
            6'd32: xpb[21] = 256'd56539106086072335005235168361013145967104442239354808069082020429944586240;
            6'd33: xpb[21] = 256'd58305953151262095474148767372294806778576456059334645821240833568380354560;
            6'd34: xpb[21] = 256'd60072800216451855943062366383576467590048469879314483573399646706816122880;
            6'd35: xpb[21] = 256'd61839647281641616411975965394858128401520483699294321325558459845251891200;
            6'd36: xpb[21] = 256'd63606494346831376880889564406139789212992497519274159077717272983687659520;
            6'd37: xpb[21] = 256'd65373341412021137349803163417421450024464511339253996829876086122123427840;
            6'd38: xpb[21] = 256'd67140188477210897818716762428703110835936525159233834582034899260559196160;
            6'd39: xpb[21] = 256'd68907035542400658287630361439984771647408538979213672334193712398994964480;
            6'd40: xpb[21] = 256'd70673882607590418756543960451266432458880552799193510086352525537430732800;
            6'd41: xpb[21] = 256'd72440729672780179225457559462548093270352566619173347838511338675866501120;
            6'd42: xpb[21] = 256'd74207576737969939694371158473829754081824580439153185590670151814302269440;
            6'd43: xpb[21] = 256'd75974423803159700163284757485111414893296594259133023342828964952738037760;
            6'd44: xpb[21] = 256'd77741270868349460632198356496393075704768608079112861094987778091173806080;
            6'd45: xpb[21] = 256'd79508117933539221101111955507674736516240621899092698847146591229609574400;
            6'd46: xpb[21] = 256'd81274964998728981570025554518956397327712635719072536599305404368045342720;
            6'd47: xpb[21] = 256'd83041812063918742038939153530238058139184649539052374351464217506481111040;
            6'd48: xpb[21] = 256'd84808659129108502507852752541519718950656663359032212103623030644916879360;
            6'd49: xpb[21] = 256'd86575506194298262976766351552801379762128677179012049855781843783352647680;
            6'd50: xpb[21] = 256'd88342353259488023445679950564083040573600690998991887607940656921788416000;
            6'd51: xpb[21] = 256'd90109200324677783914593549575364701385072704818971725360099470060224184320;
            6'd52: xpb[21] = 256'd91876047389867544383507148586646362196544718638951563112258283198659952640;
            6'd53: xpb[21] = 256'd93642894455057304852420747597928023008016732458931400864417096337095720960;
            6'd54: xpb[21] = 256'd95409741520247065321334346609209683819488746278911238616575909475531489280;
            6'd55: xpb[21] = 256'd97176588585436825790247945620491344630960760098891076368734722613967257600;
            6'd56: xpb[21] = 256'd98943435650626586259161544631773005442432773918870914120893535752403025920;
            6'd57: xpb[21] = 256'd100710282715816346728075143643054666253904787738850751873052348890838794240;
            6'd58: xpb[21] = 256'd102477129781006107196988742654336327065376801558830589625211162029274562560;
            6'd59: xpb[21] = 256'd104243976846195867665902341665617987876848815378810427377369975167710330880;
            6'd60: xpb[21] = 256'd106010823911385628134815940676899648688320829198790265129528788306146099200;
            6'd61: xpb[21] = 256'd107777670976575388603729539688181309499792843018770102881687601444581867520;
            6'd62: xpb[21] = 256'd109544518041765149072643138699462970311264856838749940633846414583017635840;
            6'd63: xpb[21] = 256'd111311365106954909541556737710744631122736870658729778386005227721453404160;
        endcase
    end

    always_comb begin
        case(flag[22])
            6'd0: xpb[22] = 256'd0;
            6'd1: xpb[22] = 256'd113078212172144670010470336722026291934208884478709616138164040859889172480;
            6'd2: xpb[22] = 256'd226156424344289340020940673444052583868417768957419232276328081719778344960;
            6'd3: xpb[22] = 256'd339234636516434010031411010166078875802626653436128848414492122579667517440;
            6'd4: xpb[22] = 256'd452312848688578680041881346888105167736835537914838464552656163439556689920;
            6'd5: xpb[22] = 256'd565391060860723350052351683610131459671044422393548080690820204299445862400;
            6'd6: xpb[22] = 256'd678469273032868020062822020332157751605253306872257696828984245159335034880;
            6'd7: xpb[22] = 256'd791547485205012690073292357054184043539462191350967312967148286019224207360;
            6'd8: xpb[22] = 256'd904625697377157360083762693776210335473671075829676929105312326879113379840;
            6'd9: xpb[22] = 256'd1017703909549302030094233030498236627407879960308386545243476367739002552320;
            6'd10: xpb[22] = 256'd1130782121721446700104703367220262919342088844787096161381640408598891724800;
            6'd11: xpb[22] = 256'd1243860333893591370115173703942289211276297729265805777519804449458780897280;
            6'd12: xpb[22] = 256'd1356938546065736040125644040664315503210506613744515393657968490318670069760;
            6'd13: xpb[22] = 256'd1470016758237880710136114377386341795144715498223225009796132531178559242240;
            6'd14: xpb[22] = 256'd1583094970410025380146584714108368087078924382701934625934296572038448414720;
            6'd15: xpb[22] = 256'd1696173182582170050157055050830394379013133267180644242072460612898337587200;
            6'd16: xpb[22] = 256'd1809251394754314720167525387552420670947342151659353858210624653758226759680;
            6'd17: xpb[22] = 256'd1922329606926459390177995724274446962881551036138063474348788694618115932160;
            6'd18: xpb[22] = 256'd2035407819098604060188466060996473254815759920616773090486952735478005104640;
            6'd19: xpb[22] = 256'd2148486031270748730198936397718499546749968805095482706625116776337894277120;
            6'd20: xpb[22] = 256'd2261564243442893400209406734440525838684177689574192322763280817197783449600;
            6'd21: xpb[22] = 256'd2374642455615038070219877071162552130618386574052901938901444858057672622080;
            6'd22: xpb[22] = 256'd2487720667787182740230347407884578422552595458531611555039608898917561794560;
            6'd23: xpb[22] = 256'd2600798879959327410240817744606604714486804343010321171177772939777450967040;
            6'd24: xpb[22] = 256'd2713877092131472080251288081328631006421013227489030787315936980637340139520;
            6'd25: xpb[22] = 256'd2826955304303616750261758418050657298355222111967740403454101021497229312000;
            6'd26: xpb[22] = 256'd2940033516475761420272228754772683590289430996446450019592265062357118484480;
            6'd27: xpb[22] = 256'd3053111728647906090282699091494709882223639880925159635730429103217007656960;
            6'd28: xpb[22] = 256'd3166189940820050760293169428216736174157848765403869251868593144076896829440;
            6'd29: xpb[22] = 256'd3279268152992195430303639764938762466092057649882578868006757184936786001920;
            6'd30: xpb[22] = 256'd3392346365164340100314110101660788758026266534361288484144921225796675174400;
            6'd31: xpb[22] = 256'd3505424577336484770324580438382815049960475418839998100283085266656564346880;
            6'd32: xpb[22] = 256'd3618502789508629440335050775104841341894684303318707716421249307516453519360;
            6'd33: xpb[22] = 256'd3731581001680774110345521111826867633828893187797417332559413348376342691840;
            6'd34: xpb[22] = 256'd3844659213852918780355991448548893925763102072276126948697577389236231864320;
            6'd35: xpb[22] = 256'd3957737426025063450366461785270920217697310956754836564835741430096121036800;
            6'd36: xpb[22] = 256'd4070815638197208120376932121992946509631519841233546180973905470956010209280;
            6'd37: xpb[22] = 256'd4183893850369352790387402458714972801565728725712255797112069511815899381760;
            6'd38: xpb[22] = 256'd4296972062541497460397872795436999093499937610190965413250233552675788554240;
            6'd39: xpb[22] = 256'd4410050274713642130408343132159025385434146494669675029388397593535677726720;
            6'd40: xpb[22] = 256'd4523128486885786800418813468881051677368355379148384645526561634395566899200;
            6'd41: xpb[22] = 256'd4636206699057931470429283805603077969302564263627094261664725675255456071680;
            6'd42: xpb[22] = 256'd4749284911230076140439754142325104261236773148105803877802889716115345244160;
            6'd43: xpb[22] = 256'd4862363123402220810450224479047130553170982032584513493941053756975234416640;
            6'd44: xpb[22] = 256'd4975441335574365480460694815769156845105190917063223110079217797835123589120;
            6'd45: xpb[22] = 256'd5088519547746510150471165152491183137039399801541932726217381838695012761600;
            6'd46: xpb[22] = 256'd5201597759918654820481635489213209428973608686020642342355545879554901934080;
            6'd47: xpb[22] = 256'd5314675972090799490492105825935235720907817570499351958493709920414791106560;
            6'd48: xpb[22] = 256'd5427754184262944160502576162657262012842026454978061574631873961274680279040;
            6'd49: xpb[22] = 256'd5540832396435088830513046499379288304776235339456771190770038002134569451520;
            6'd50: xpb[22] = 256'd5653910608607233500523516836101314596710444223935480806908202042994458624000;
            6'd51: xpb[22] = 256'd5766988820779378170533987172823340888644653108414190423046366083854347796480;
            6'd52: xpb[22] = 256'd5880067032951522840544457509545367180578861992892900039184530124714236968960;
            6'd53: xpb[22] = 256'd5993145245123667510554927846267393472513070877371609655322694165574126141440;
            6'd54: xpb[22] = 256'd6106223457295812180565398182989419764447279761850319271460858206434015313920;
            6'd55: xpb[22] = 256'd6219301669467956850575868519711446056381488646329028887599022247293904486400;
            6'd56: xpb[22] = 256'd6332379881640101520586338856433472348315697530807738503737186288153793658880;
            6'd57: xpb[22] = 256'd6445458093812246190596809193155498640249906415286448119875350329013682831360;
            6'd58: xpb[22] = 256'd6558536305984390860607279529877524932184115299765157736013514369873572003840;
            6'd59: xpb[22] = 256'd6671614518156535530617749866599551224118324184243867352151678410733461176320;
            6'd60: xpb[22] = 256'd6784692730328680200628220203321577516052533068722576968289842451593350348800;
            6'd61: xpb[22] = 256'd6897770942500824870638690540043603807986741953201286584428006492453239521280;
            6'd62: xpb[22] = 256'd7010849154672969540649160876765630099920950837679996200566170533313128693760;
            6'd63: xpb[22] = 256'd7123927366845114210659631213487656391855159722158705816704334574173017866240;
        endcase
    end

    always_comb begin
        case(flag[23])
            6'd0: xpb[23] = 256'd0;
            6'd1: xpb[23] = 256'd7237005579017258880670101550209682683789368606637415432842498615032907038720;
            6'd2: xpb[23] = 256'd14474011158034517761340203100419365367578737213274830865684997230065814077440;
            6'd3: xpb[23] = 256'd21711016737051776642010304650629048051368105819912246298527495845098721116160;
            6'd4: xpb[23] = 256'd28948022316069035522680406200838730735157474426549661731369994460131628154880;
            6'd5: xpb[23] = 256'd36185027895086294403350507751048413418946843033187077164212493075164535193600;
            6'd6: xpb[23] = 256'd43422033474103553284020609301258096102736211639824492597054991690197442232320;
            6'd7: xpb[23] = 256'd50659039053120812164690710851467778786525580246461908029897490305230349271040;
            6'd8: xpb[23] = 256'd57896044632138071045360812401677461470314948853099323462739988920263256309760;
            6'd9: xpb[23] = 256'd65133050211155329926030913951887144154104317459736738895582487535296163348480;
            6'd10: xpb[23] = 256'd72370055790172588806701015502096826837893686066374154328424986150329070387200;
            6'd11: xpb[23] = 256'd79607061369189847687371117052306509521683054673011569761267484765361977425920;
            6'd12: xpb[23] = 256'd86844066948207106568041218602516192205472423279648985194109983380394884464640;
            6'd13: xpb[23] = 256'd94081072527224365448711320152725874889261791886286400626952481995427791503360;
            6'd14: xpb[23] = 256'd101318078106241624329381421702935557573051160492923816059794980610460698542080;
            6'd15: xpb[23] = 256'd108555083685258883210051523253145240256840529099561231492637479225493605580800;
            6'd16: xpb[23] = 256'd53919893334301279589334030174379543714274455471058783907236827627521;
            6'd17: xpb[23] = 256'd7237005632937152214971381139543712858168912320911870903901282522269734666241;
            6'd18: xpb[23] = 256'd14474011211954411095641482689753395541958280927549286336743781137302641704961;
            6'd19: xpb[23] = 256'd21711016790971669976311584239963078225747649534186701769586279752335548743681;
            6'd20: xpb[23] = 256'd28948022369988928856981685790172760909537018140824117202428778367368455782401;
            6'd21: xpb[23] = 256'd36185027949006187737651787340382443593326386747461532635271276982401362821121;
            6'd22: xpb[23] = 256'd43422033528023446618321888890592126277115755354098948068113775597434269859841;
            6'd23: xpb[23] = 256'd50659039107040705498991990440801808960905123960736363500956274212467176898561;
            6'd24: xpb[23] = 256'd57896044686057964379662091991011491644694492567373778933798772827500083937281;
            6'd25: xpb[23] = 256'd65133050265075223260332193541221174328483861174011194366641271442532990976001;
            6'd26: xpb[23] = 256'd72370055844092482141002295091430857012273229780648609799483770057565898014721;
            6'd27: xpb[23] = 256'd79607061423109741021672396641640539696062598387286025232326268672598805053441;
            6'd28: xpb[23] = 256'd86844067002126999902342498191850222379851966993923440665168767287631712092161;
            6'd29: xpb[23] = 256'd94081072581144258783012599742059905063641335600560856098011265902664619130881;
            6'd30: xpb[23] = 256'd101318078160161517663682701292269587747430704207198271530853764517697526169601;
            6'd31: xpb[23] = 256'd108555083739178776544352802842479270431220072813835686963696263132730433208321;
            6'd32: xpb[23] = 256'd107839786668602559178668060348759087428548910942117567814473655255042;
            6'd33: xpb[23] = 256'd7237005686857045549272660728877743032548456035186326374960066429506562293762;
            6'd34: xpb[23] = 256'd14474011265874304429942762279087425716337824641823741807802565044539469332482;
            6'd35: xpb[23] = 256'd21711016844891563310612863829297108400127193248461157240645063659572376371202;
            6'd36: xpb[23] = 256'd28948022423908822191282965379506791083916561855098572673487562274605283409922;
            6'd37: xpb[23] = 256'd36185028002926081071953066929716473767705930461735988106330060889638190448642;
            6'd38: xpb[23] = 256'd43422033581943339952623168479926156451495299068373403539172559504671097487362;
            6'd39: xpb[23] = 256'd50659039160960598833293270030135839135284667675010818972015058119704004526082;
            6'd40: xpb[23] = 256'd57896044739977857713963371580345521819074036281648234404857556734736911564802;
            6'd41: xpb[23] = 256'd65133050318995116594633473130555204502863404888285649837700055349769818603522;
            6'd42: xpb[23] = 256'd72370055898012375475303574680764887186652773494923065270542553964802725642242;
            6'd43: xpb[23] = 256'd79607061477029634355973676230974569870442142101560480703385052579835632680962;
            6'd44: xpb[23] = 256'd86844067056046893236643777781184252554231510708197896136227551194868539719682;
            6'd45: xpb[23] = 256'd94081072635064152117313879331393935238020879314835311569070049809901446758402;
            6'd46: xpb[23] = 256'd101318078214081410997983980881603617921810247921472727001912548424934353797122;
            6'd47: xpb[23] = 256'd108555083793098669878654082431813300605599616528110142434755047039967260835842;
            6'd48: xpb[23] = 256'd161759680002903838768002090523138631142823366413176351721710482882563;
            6'd49: xpb[23] = 256'd7237005740776938883573940318211773206927999749460781846018850336743389921283;
            6'd50: xpb[23] = 256'd14474011319794197764244041868421455890717368356098197278861348951776296960003;
            6'd51: xpb[23] = 256'd21711016898811456644914143418631138574506736962735612711703847566809203998723;
            6'd52: xpb[23] = 256'd28948022477828715525584244968840821258296105569373028144546346181842111037443;
            6'd53: xpb[23] = 256'd36185028056845974406254346519050503942085474176010443577388844796875018076163;
            6'd54: xpb[23] = 256'd43422033635863233286924448069260186625874842782647859010231343411907925114883;
            6'd55: xpb[23] = 256'd50659039214880492167594549619469869309664211389285274443073842026940832153603;
            6'd56: xpb[23] = 256'd57896044793897751048264651169679551993453579995922689875916340641973739192323;
            6'd57: xpb[23] = 256'd65133050372915009928934752719889234677242948602560105308758839257006646231043;
            6'd58: xpb[23] = 256'd72370055951932268809604854270098917361032317209197520741601337872039553269763;
            6'd59: xpb[23] = 256'd79607061530949527690274955820308600044821685815834936174443836487072460308483;
            6'd60: xpb[23] = 256'd86844067109966786570945057370518282728611054422472351607286335102105367347203;
            6'd61: xpb[23] = 256'd94081072688984045451615158920727965412400423029109767040128833717138274385923;
            6'd62: xpb[23] = 256'd101318078268001304332285260470937648096189791635747182472971332332171181424643;
            6'd63: xpb[23] = 256'd108555083847018563212955362021147330779979160242384597905813830947204088463363;
        endcase
    end

    always_comb begin
        case(flag[24])
            6'd0: xpb[24] = 256'd0;
            6'd1: xpb[24] = 256'd53919893334301279589334030174379543714274455471058783907236827627521;
            6'd2: xpb[24] = 256'd107839786668602559178668060348759087428548910942117567814473655255042;
            6'd3: xpb[24] = 256'd161759680002903838768002090523138631142823366413176351721710482882563;
            6'd4: xpb[24] = 256'd215679573337205118357336120697518174857097821884235135628947310510084;
            6'd5: xpb[24] = 256'd269599466671506397946670150871897718571372277355293919536184138137605;
            6'd6: xpb[24] = 256'd323519360005807677536004181046277262285646732826352703443420965765126;
            6'd7: xpb[24] = 256'd377439253340108957125338211220656805999921188297411487350657793392647;
            6'd8: xpb[24] = 256'd431359146674410236714672241395036349714195643768470271257894621020168;
            6'd9: xpb[24] = 256'd485279040008711516304006271569415893428470099239529055165131448647689;
            6'd10: xpb[24] = 256'd539198933343012795893340301743795437142744554710587839072368276275210;
            6'd11: xpb[24] = 256'd593118826677314075482674331918174980857019010181646622979605103902731;
            6'd12: xpb[24] = 256'd647038720011615355072008362092554524571293465652705406886841931530252;
            6'd13: xpb[24] = 256'd700958613345916634661342392266934068285567921123764190794078759157773;
            6'd14: xpb[24] = 256'd754878506680217914250676422441313611999842376594822974701315586785294;
            6'd15: xpb[24] = 256'd808798400014519193840010452615693155714116832065881758608552414412815;
            6'd16: xpb[24] = 256'd862718293348820473429344482790072699428391287536940542515789242040336;
            6'd17: xpb[24] = 256'd916638186683121753018678512964452243142665743007999326423026069667857;
            6'd18: xpb[24] = 256'd970558080017423032608012543138831786856940198479058110330262897295378;
            6'd19: xpb[24] = 256'd1024477973351724312197346573313211330571214653950116894237499724922899;
            6'd20: xpb[24] = 256'd1078397866686025591786680603487590874285489109421175678144736552550420;
            6'd21: xpb[24] = 256'd1132317760020326871376014633661970417999763564892234462051973380177941;
            6'd22: xpb[24] = 256'd1186237653354628150965348663836349961714038020363293245959210207805462;
            6'd23: xpb[24] = 256'd1240157546688929430554682694010729505428312475834352029866447035432983;
            6'd24: xpb[24] = 256'd1294077440023230710144016724185109049142586931305410813773683863060504;
            6'd25: xpb[24] = 256'd1347997333357531989733350754359488592856861386776469597680920690688025;
            6'd26: xpb[24] = 256'd1401917226691833269322684784533868136571135842247528381588157518315546;
            6'd27: xpb[24] = 256'd1455837120026134548912018814708247680285410297718587165495394345943067;
            6'd28: xpb[24] = 256'd1509757013360435828501352844882627223999684753189645949402631173570588;
            6'd29: xpb[24] = 256'd1563676906694737108090686875057006767713959208660704733309868001198109;
            6'd30: xpb[24] = 256'd1617596800029038387680020905231386311428233664131763517217104828825630;
            6'd31: xpb[24] = 256'd1671516693363339667269354935405765855142508119602822301124341656453151;
            6'd32: xpb[24] = 256'd1725436586697640946858688965580145398856782575073881085031578484080672;
            6'd33: xpb[24] = 256'd1779356480031942226448022995754524942571057030544939868938815311708193;
            6'd34: xpb[24] = 256'd1833276373366243506037357025928904486285331486015998652846052139335714;
            6'd35: xpb[24] = 256'd1887196266700544785626691056103284029999605941487057436753288966963235;
            6'd36: xpb[24] = 256'd1941116160034846065216025086277663573713880396958116220660525794590756;
            6'd37: xpb[24] = 256'd1995036053369147344805359116452043117428154852429175004567762622218277;
            6'd38: xpb[24] = 256'd2048955946703448624394693146626422661142429307900233788474999449845798;
            6'd39: xpb[24] = 256'd2102875840037749903984027176800802204856703763371292572382236277473319;
            6'd40: xpb[24] = 256'd2156795733372051183573361206975181748570978218842351356289473105100840;
            6'd41: xpb[24] = 256'd2210715626706352463162695237149561292285252674313410140196709932728361;
            6'd42: xpb[24] = 256'd2264635520040653742752029267323940835999527129784468924103946760355882;
            6'd43: xpb[24] = 256'd2318555413374955022341363297498320379713801585255527708011183587983403;
            6'd44: xpb[24] = 256'd2372475306709256301930697327672699923428076040726586491918420415610924;
            6'd45: xpb[24] = 256'd2426395200043557581520031357847079467142350496197645275825657243238445;
            6'd46: xpb[24] = 256'd2480315093377858861109365388021459010856624951668704059732894070865966;
            6'd47: xpb[24] = 256'd2534234986712160140698699418195838554570899407139762843640130898493487;
            6'd48: xpb[24] = 256'd2588154880046461420288033448370218098285173862610821627547367726121008;
            6'd49: xpb[24] = 256'd2642074773380762699877367478544597641999448318081880411454604553748529;
            6'd50: xpb[24] = 256'd2695994666715063979466701508718977185713722773552939195361841381376050;
            6'd51: xpb[24] = 256'd2749914560049365259056035538893356729427997229023997979269078209003571;
            6'd52: xpb[24] = 256'd2803834453383666538645369569067736273142271684495056763176315036631092;
            6'd53: xpb[24] = 256'd2857754346717967818234703599242115816856546139966115547083551864258613;
            6'd54: xpb[24] = 256'd2911674240052269097824037629416495360570820595437174330990788691886134;
            6'd55: xpb[24] = 256'd2965594133386570377413371659590874904285095050908233114898025519513655;
            6'd56: xpb[24] = 256'd3019514026720871657002705689765254447999369506379291898805262347141176;
            6'd57: xpb[24] = 256'd3073433920055172936592039719939633991713643961850350682712499174768697;
            6'd58: xpb[24] = 256'd3127353813389474216181373750114013535427918417321409466619736002396218;
            6'd59: xpb[24] = 256'd3181273706723775495770707780288393079142192872792468250526972830023739;
            6'd60: xpb[24] = 256'd3235193600058076775360041810462772622856467328263527034434209657651260;
            6'd61: xpb[24] = 256'd3289113493392378054949375840637152166570741783734585818341446485278781;
            6'd62: xpb[24] = 256'd3343033386726679334538709870811531710285016239205644602248683312906302;
            6'd63: xpb[24] = 256'd3396953280060980614128043900985911253999290694676703386155920140533823;
        endcase
    end

    always_comb begin
        case(flag[25])
            6'd0: xpb[25] = 256'd0;
            6'd1: xpb[25] = 256'd3450873173395281893717377931160290797713565150147762170063156968161344;
            6'd2: xpb[25] = 256'd6901746346790563787434755862320581595427130300295524340126313936322688;
            6'd3: xpb[25] = 256'd10352619520185845681152133793480872393140695450443286510189470904484032;
            6'd4: xpb[25] = 256'd13803492693581127574869511724641163190854260600591048680252627872645376;
            6'd5: xpb[25] = 256'd17254365866976409468586889655801453988567825750738810850315784840806720;
            6'd6: xpb[25] = 256'd20705239040371691362304267586961744786281390900886573020378941808968064;
            6'd7: xpb[25] = 256'd24156112213766973256021645518122035583994956051034335190442098777129408;
            6'd8: xpb[25] = 256'd27606985387162255149739023449282326381708521201182097360505255745290752;
            6'd9: xpb[25] = 256'd31057858560557537043456401380442617179422086351329859530568412713452096;
            6'd10: xpb[25] = 256'd34508731733952818937173779311602907977135651501477621700631569681613440;
            6'd11: xpb[25] = 256'd37959604907348100830891157242763198774849216651625383870694726649774784;
            6'd12: xpb[25] = 256'd41410478080743382724608535173923489572562781801773146040757883617936128;
            6'd13: xpb[25] = 256'd44861351254138664618325913105083780370276346951920908210821040586097472;
            6'd14: xpb[25] = 256'd48312224427533946512043291036244071167989912102068670380884197554258816;
            6'd15: xpb[25] = 256'd51763097600929228405760668967404361965703477252216432550947354522420160;
            6'd16: xpb[25] = 256'd55213970774324510299478046898564652763417042402364194721010511490581504;
            6'd17: xpb[25] = 256'd58664843947719792193195424829724943561130607552511956891073668458742848;
            6'd18: xpb[25] = 256'd62115717121115074086912802760885234358844172702659719061136825426904192;
            6'd19: xpb[25] = 256'd65566590294510355980630180692045525156557737852807481231199982395065536;
            6'd20: xpb[25] = 256'd69017463467905637874347558623205815954271303002955243401263139363226880;
            6'd21: xpb[25] = 256'd72468336641300919768064936554366106751984868153103005571326296331388224;
            6'd22: xpb[25] = 256'd75919209814696201661782314485526397549698433303250767741389453299549568;
            6'd23: xpb[25] = 256'd79370082988091483555499692416686688347411998453398529911452610267710912;
            6'd24: xpb[25] = 256'd82820956161486765449217070347846979145125563603546292081515767235872256;
            6'd25: xpb[25] = 256'd86271829334882047342934448279007269942839128753694054251578924204033600;
            6'd26: xpb[25] = 256'd89722702508277329236651826210167560740552693903841816421642081172194944;
            6'd27: xpb[25] = 256'd93173575681672611130369204141327851538266259053989578591705238140356288;
            6'd28: xpb[25] = 256'd96624448855067893024086582072488142335979824204137340761768395108517632;
            6'd29: xpb[25] = 256'd100075322028463174917803960003648433133693389354285102931831552076678976;
            6'd30: xpb[25] = 256'd103526195201858456811521337934808723931406954504432865101894709044840320;
            6'd31: xpb[25] = 256'd106977068375253738705238715865969014729120519654580627271957866013001664;
            6'd32: xpb[25] = 256'd110427941548649020598956093797129305526834084804728389442021022981163008;
            6'd33: xpb[25] = 256'd113878814722044302492673471728289596324547649954876151612084179949324352;
            6'd34: xpb[25] = 256'd117329687895439584386390849659449887122261215105023913782147336917485696;
            6'd35: xpb[25] = 256'd120780561068834866280108227590610177919974780255171675952210493885647040;
            6'd36: xpb[25] = 256'd124231434242230148173825605521770468717688345405319438122273650853808384;
            6'd37: xpb[25] = 256'd127682307415625430067542983452930759515401910555467200292336807821969728;
            6'd38: xpb[25] = 256'd131133180589020711961260361384091050313115475705614962462399964790131072;
            6'd39: xpb[25] = 256'd134584053762415993854977739315251341110829040855762724632463121758292416;
            6'd40: xpb[25] = 256'd138034926935811275748695117246411631908542606005910486802526278726453760;
            6'd41: xpb[25] = 256'd141485800109206557642412495177571922706256171156058248972589435694615104;
            6'd42: xpb[25] = 256'd144936673282601839536129873108732213503969736306206011142652592662776448;
            6'd43: xpb[25] = 256'd148387546455997121429847251039892504301683301456353773312715749630937792;
            6'd44: xpb[25] = 256'd151838419629392403323564628971052795099396866606501535482778906599099136;
            6'd45: xpb[25] = 256'd155289292802787685217282006902213085897110431756649297652842063567260480;
            6'd46: xpb[25] = 256'd158740165976182967110999384833373376694823996906797059822905220535421824;
            6'd47: xpb[25] = 256'd162191039149578249004716762764533667492537562056944821992968377503583168;
            6'd48: xpb[25] = 256'd165641912322973530898434140695693958290251127207092584163031534471744512;
            6'd49: xpb[25] = 256'd169092785496368812792151518626854249087964692357240346333094691439905856;
            6'd50: xpb[25] = 256'd172543658669764094685868896558014539885678257507388108503157848408067200;
            6'd51: xpb[25] = 256'd175994531843159376579586274489174830683391822657535870673221005376228544;
            6'd52: xpb[25] = 256'd179445405016554658473303652420335121481105387807683632843284162344389888;
            6'd53: xpb[25] = 256'd182896278189949940367021030351495412278818952957831395013347319312551232;
            6'd54: xpb[25] = 256'd186347151363345222260738408282655703076532518107979157183410476280712576;
            6'd55: xpb[25] = 256'd189798024536740504154455786213815993874246083258126919353473633248873920;
            6'd56: xpb[25] = 256'd193248897710135786048173164144976284671959648408274681523536790217035264;
            6'd57: xpb[25] = 256'd196699770883531067941890542076136575469673213558422443693599947185196608;
            6'd58: xpb[25] = 256'd200150644056926349835607920007296866267386778708570205863663104153357952;
            6'd59: xpb[25] = 256'd203601517230321631729325297938457157065100343858717968033726261121519296;
            6'd60: xpb[25] = 256'd207052390403716913623042675869617447862813909008865730203789418089680640;
            6'd61: xpb[25] = 256'd210503263577112195516760053800777738660527474159013492373852575057841984;
            6'd62: xpb[25] = 256'd213954136750507477410477431731938029458241039309161254543915732026003328;
            6'd63: xpb[25] = 256'd217405009923902759304194809663098320255954604459309016713978888994164672;
        endcase
    end

    always_comb begin
        case(flag[26])
            6'd0: xpb[26] = 256'd0;
            6'd1: xpb[26] = 256'd220855883097298041197912187594258611053668169609456778884042045962326016;
            6'd2: xpb[26] = 256'd441711766194596082395824375188517222107336339218913557768084091924652032;
            6'd3: xpb[26] = 256'd662567649291894123593736562782775833161004508828370336652126137886978048;
            6'd4: xpb[26] = 256'd883423532389192164791648750377034444214672678437827115536168183849304064;
            6'd5: xpb[26] = 256'd1104279415486490205989560937971293055268340848047283894420210229811630080;
            6'd6: xpb[26] = 256'd1325135298583788247187473125565551666322009017656740673304252275773956096;
            6'd7: xpb[26] = 256'd1545991181681086288385385313159810277375677187266197452188294321736282112;
            6'd8: xpb[26] = 256'd1766847064778384329583297500754068888429345356875654231072336367698608128;
            6'd9: xpb[26] = 256'd1987702947875682370781209688348327499483013526485111009956378413660934144;
            6'd10: xpb[26] = 256'd2208558830972980411979121875942586110536681696094567788840420459623260160;
            6'd11: xpb[26] = 256'd2429414714070278453177034063536844721590349865704024567724462505585586176;
            6'd12: xpb[26] = 256'd2650270597167576494374946251131103332644018035313481346608504551547912192;
            6'd13: xpb[26] = 256'd2871126480264874535572858438725361943697686204922938125492546597510238208;
            6'd14: xpb[26] = 256'd3091982363362172576770770626319620554751354374532394904376588643472564224;
            6'd15: xpb[26] = 256'd3312838246459470617968682813913879165805022544141851683260630689434890240;
            6'd16: xpb[26] = 256'd3533694129556768659166595001508137776858690713751308462144672735397216256;
            6'd17: xpb[26] = 256'd3754550012654066700364507189102396387912358883360765241028714781359542272;
            6'd18: xpb[26] = 256'd3975405895751364741562419376696654998966027052970222019912756827321868288;
            6'd19: xpb[26] = 256'd4196261778848662782760331564290913610019695222579678798796798873284194304;
            6'd20: xpb[26] = 256'd4417117661945960823958243751885172221073363392189135577680840919246520320;
            6'd21: xpb[26] = 256'd4637973545043258865156155939479430832127031561798592356564882965208846336;
            6'd22: xpb[26] = 256'd4858829428140556906354068127073689443180699731408049135448925011171172352;
            6'd23: xpb[26] = 256'd5079685311237854947551980314667948054234367901017505914332967057133498368;
            6'd24: xpb[26] = 256'd5300541194335152988749892502262206665288036070626962693217009103095824384;
            6'd25: xpb[26] = 256'd5521397077432451029947804689856465276341704240236419472101051149058150400;
            6'd26: xpb[26] = 256'd5742252960529749071145716877450723887395372409845876250985093195020476416;
            6'd27: xpb[26] = 256'd5963108843627047112343629065044982498449040579455333029869135240982802432;
            6'd28: xpb[26] = 256'd6183964726724345153541541252639241109502708749064789808753177286945128448;
            6'd29: xpb[26] = 256'd6404820609821643194739453440233499720556376918674246587637219332907454464;
            6'd30: xpb[26] = 256'd6625676492918941235937365627827758331610045088283703366521261378869780480;
            6'd31: xpb[26] = 256'd6846532376016239277135277815422016942663713257893160145405303424832106496;
            6'd32: xpb[26] = 256'd7067388259113537318333190003016275553717381427502616924289345470794432512;
            6'd33: xpb[26] = 256'd7288244142210835359531102190610534164771049597112073703173387516756758528;
            6'd34: xpb[26] = 256'd7509100025308133400729014378204792775824717766721530482057429562719084544;
            6'd35: xpb[26] = 256'd7729955908405431441926926565799051386878385936330987260941471608681410560;
            6'd36: xpb[26] = 256'd7950811791502729483124838753393309997932054105940444039825513654643736576;
            6'd37: xpb[26] = 256'd8171667674600027524322750940987568608985722275549900818709555700606062592;
            6'd38: xpb[26] = 256'd8392523557697325565520663128581827220039390445159357597593597746568388608;
            6'd39: xpb[26] = 256'd8613379440794623606718575316176085831093058614768814376477639792530714624;
            6'd40: xpb[26] = 256'd8834235323891921647916487503770344442146726784378271155361681838493040640;
            6'd41: xpb[26] = 256'd9055091206989219689114399691364603053200394953987727934245723884455366656;
            6'd42: xpb[26] = 256'd9275947090086517730312311878958861664254063123597184713129765930417692672;
            6'd43: xpb[26] = 256'd9496802973183815771510224066553120275307731293206641492013807976380018688;
            6'd44: xpb[26] = 256'd9717658856281113812708136254147378886361399462816098270897850022342344704;
            6'd45: xpb[26] = 256'd9938514739378411853906048441741637497415067632425555049781892068304670720;
            6'd46: xpb[26] = 256'd10159370622475709895103960629335896108468735802035011828665934114266996736;
            6'd47: xpb[26] = 256'd10380226505573007936301872816930154719522403971644468607549976160229322752;
            6'd48: xpb[26] = 256'd10601082388670305977499785004524413330576072141253925386434018206191648768;
            6'd49: xpb[26] = 256'd10821938271767604018697697192118671941629740310863382165318060252153974784;
            6'd50: xpb[26] = 256'd11042794154864902059895609379712930552683408480472838944202102298116300800;
            6'd51: xpb[26] = 256'd11263650037962200101093521567307189163737076650082295723086144344078626816;
            6'd52: xpb[26] = 256'd11484505921059498142291433754901447774790744819691752501970186390040952832;
            6'd53: xpb[26] = 256'd11705361804156796183489345942495706385844412989301209280854228436003278848;
            6'd54: xpb[26] = 256'd11926217687254094224687258130089964996898081158910666059738270481965604864;
            6'd55: xpb[26] = 256'd12147073570351392265885170317684223607951749328520122838622312527927930880;
            6'd56: xpb[26] = 256'd12367929453448690307083082505278482219005417498129579617506354573890256896;
            6'd57: xpb[26] = 256'd12588785336545988348280994692872740830059085667739036396390396619852582912;
            6'd58: xpb[26] = 256'd12809641219643286389478906880466999441112753837348493175274438665814908928;
            6'd59: xpb[26] = 256'd13030497102740584430676819068061258052166422006957949954158480711777234944;
            6'd60: xpb[26] = 256'd13251352985837882471874731255655516663220090176567406733042522757739560960;
            6'd61: xpb[26] = 256'd13472208868935180513072643443249775274273758346176863511926564803701886976;
            6'd62: xpb[26] = 256'd13693064752032478554270555630844033885327426515786320290810606849664212992;
            6'd63: xpb[26] = 256'd13913920635129776595468467818438292496381094685395777069694648895626539008;
        endcase
    end

    always_comb begin
        case(flag[27])
            6'd0: xpb[27] = 256'd0;
            6'd1: xpb[27] = 256'd3533694129556768659166595001508137776858690713751308462144672735397216256;
            6'd2: xpb[27] = 256'd7067388259113537318333190003016275553717381427502616924289345470794432512;
            6'd3: xpb[27] = 256'd10601082388670305977499785004524413330576072141253925386434018206191648768;
            6'd4: xpb[27] = 256'd14134776518227074636666380006032551107434762855005233848578690941588865024;
            6'd5: xpb[27] = 256'd17668470647783843295832975007540688884293453568756542310723363676986081280;
            6'd6: xpb[27] = 256'd21202164777340611954999570009048826661152144282507850772868036412383297536;
            6'd7: xpb[27] = 256'd24735858906897380614166165010556964438010834996259159235012709147780513792;
            6'd8: xpb[27] = 256'd28269553036454149273332760012065102214869525710010467697157381883177730048;
            6'd9: xpb[27] = 256'd31803247166010917932499355013573239991728216423761776159302054618574946304;
            6'd10: xpb[27] = 256'd35336941295567686591665950015081377768586907137513084621446727353972162560;
            6'd11: xpb[27] = 256'd38870635425124455250832545016589515545445597851264393083591400089369378816;
            6'd12: xpb[27] = 256'd42404329554681223909999140018097653322304288565015701545736072824766595072;
            6'd13: xpb[27] = 256'd45938023684237992569165735019605791099162979278767010007880745560163811328;
            6'd14: xpb[27] = 256'd49471717813794761228332330021113928876021669992518318470025418295561027584;
            6'd15: xpb[27] = 256'd53005411943351529887498925022622066652880360706269626932170091030958243840;
            6'd16: xpb[27] = 256'd56539106072908298546665520024130204429739051420020935394314763766355460096;
            6'd17: xpb[27] = 256'd60072800202465067205832115025638342206597742133772243856459436501752676352;
            6'd18: xpb[27] = 256'd63606494332021835864998710027146479983456432847523552318604109237149892608;
            6'd19: xpb[27] = 256'd67140188461578604524165305028654617760315123561274860780748781972547108864;
            6'd20: xpb[27] = 256'd70673882591135373183331900030162755537173814275026169242893454707944325120;
            6'd21: xpb[27] = 256'd74207576720692141842498495031670893314032504988777477705038127443341541376;
            6'd22: xpb[27] = 256'd77741270850248910501665090033179031090891195702528786167182800178738757632;
            6'd23: xpb[27] = 256'd81274964979805679160831685034687168867749886416280094629327472914135973888;
            6'd24: xpb[27] = 256'd84808659109362447819998280036195306644608577130031403091472145649533190144;
            6'd25: xpb[27] = 256'd88342353238919216479164875037703444421467267843782711553616818384930406400;
            6'd26: xpb[27] = 256'd91876047368475985138331470039211582198325958557534020015761491120327622656;
            6'd27: xpb[27] = 256'd95409741498032753797498065040719719975184649271285328477906163855724838912;
            6'd28: xpb[27] = 256'd98943435627589522456664660042227857752043339985036636940050836591122055168;
            6'd29: xpb[27] = 256'd102477129757146291115831255043735995528902030698787945402195509326519271424;
            6'd30: xpb[27] = 256'd106010823886703059774997850045244133305760721412539253864340182061916487680;
            6'd31: xpb[27] = 256'd109544518016259828434164445046752271082619412126290562326484854797313703936;
            6'd32: xpb[27] = 256'd113078212145816597093331040048260408859478102840041870788629527532710920192;
            6'd33: xpb[27] = 256'd116611906275373365752497635049768546636336793553793179250774200268108136448;
            6'd34: xpb[27] = 256'd120145600404930134411664230051276684413195484267544487712918873003505352704;
            6'd35: xpb[27] = 256'd123679294534486903070830825052784822190054174981295796175063545738902568960;
            6'd36: xpb[27] = 256'd127212988664043671729997420054292959966912865695047104637208218474299785216;
            6'd37: xpb[27] = 256'd130746682793600440389164015055801097743771556408798413099352891209697001472;
            6'd38: xpb[27] = 256'd134280376923157209048330610057309235520630247122549721561497563945094217728;
            6'd39: xpb[27] = 256'd137814071052713977707497205058817373297488937836301030023642236680491433984;
            6'd40: xpb[27] = 256'd141347765182270746366663800060325511074347628550052338485786909415888650240;
            6'd41: xpb[27] = 256'd144881459311827515025830395061833648851206319263803646947931582151285866496;
            6'd42: xpb[27] = 256'd148415153441384283684996990063341786628065009977554955410076254886683082752;
            6'd43: xpb[27] = 256'd151948847570941052344163585064849924404923700691306263872220927622080299008;
            6'd44: xpb[27] = 256'd155482541700497821003330180066358062181782391405057572334365600357477515264;
            6'd45: xpb[27] = 256'd159016235830054589662496775067866199958641082118808880796510273092874731520;
            6'd46: xpb[27] = 256'd162549929959611358321663370069374337735499772832560189258654945828271947776;
            6'd47: xpb[27] = 256'd166083624089168126980829965070882475512358463546311497720799618563669164032;
            6'd48: xpb[27] = 256'd169617318218724895639996560072390613289217154260062806182944291299066380288;
            6'd49: xpb[27] = 256'd173151012348281664299163155073898751066075844973814114645088964034463596544;
            6'd50: xpb[27] = 256'd176684706477838432958329750075406888842934535687565423107233636769860812800;
            6'd51: xpb[27] = 256'd180218400607395201617496345076915026619793226401316731569378309505258029056;
            6'd52: xpb[27] = 256'd183752094736951970276662940078423164396651917115068040031522982240655245312;
            6'd53: xpb[27] = 256'd187285788866508738935829535079931302173510607828819348493667654976052461568;
            6'd54: xpb[27] = 256'd190819482996065507594996130081439439950369298542570656955812327711449677824;
            6'd55: xpb[27] = 256'd194353177125622276254162725082947577727227989256321965417957000446846894080;
            6'd56: xpb[27] = 256'd197886871255179044913329320084455715504086679970073273880101673182244110336;
            6'd57: xpb[27] = 256'd201420565384735813572495915085963853280945370683824582342246345917641326592;
            6'd58: xpb[27] = 256'd204954259514292582231662510087471991057804061397575890804391018653038542848;
            6'd59: xpb[27] = 256'd208487953643849350890829105088980128834662752111327199266535691388435759104;
            6'd60: xpb[27] = 256'd212021647773406119549995700090488266611521442825078507728680364123832975360;
            6'd61: xpb[27] = 256'd215555341902962888209162295091996404388380133538829816190825036859230191616;
            6'd62: xpb[27] = 256'd219089036032519656868328890093504542165238824252581124652969709594627407872;
            6'd63: xpb[27] = 256'd222622730162076425527495485095012679942097514966332433115114382330024624128;
        endcase
    end

    always_comb begin
        case(flag[28])
            6'd0: xpb[28] = 256'd0;
            6'd1: xpb[28] = 256'd226156424291633194186662080096520817718956205680083741577259055065421840384;
            6'd2: xpb[28] = 256'd452312848583266388373324160193041635437912411360167483154518110130843680768;
            6'd3: xpb[28] = 256'd678469272874899582559986240289562453156868617040251224731777165196265521152;
            6'd4: xpb[28] = 256'd904625697166532776746648320386083270875824822720334966309036220261687361536;
            6'd5: xpb[28] = 256'd1130782121458165970933310400482604088594781028400418707886295275327109201920;
            6'd6: xpb[28] = 256'd1356938545749799165119972480579124906313737234080502449463554330392531042304;
            6'd7: xpb[28] = 256'd1583094970041432359306634560675645724032693439760586191040813385457952882688;
            6'd8: xpb[28] = 256'd1809251394333065553493296640772166541751649645440669932618072440523374723072;
            6'd9: xpb[28] = 256'd2035407818624698747679958720868687359470605851120753674195331495588796563456;
            6'd10: xpb[28] = 256'd2261564242916331941866620800965208177189562056800837415772590550654218403840;
            6'd11: xpb[28] = 256'd2487720667207965136053282881061728994908518262480921157349849605719640244224;
            6'd12: xpb[28] = 256'd2713877091499598330239944961158249812627474468161004898927108660785062084608;
            6'd13: xpb[28] = 256'd2940033515791231524426607041254770630346430673841088640504367715850483924992;
            6'd14: xpb[28] = 256'd3166189940082864718613269121351291448065386879521172382081626770915905765376;
            6'd15: xpb[28] = 256'd3392346364374497912799931201447812265784343085201256123658885825981327605760;
            6'd16: xpb[28] = 256'd3618502788666131106986593281544333083503299290881339865236144881046749446144;
            6'd17: xpb[28] = 256'd3844659212957764301173255361640853901222255496561423606813403936112171286528;
            6'd18: xpb[28] = 256'd4070815637249397495359917441737374718941211702241507348390662991177593126912;
            6'd19: xpb[28] = 256'd4296972061541030689546579521833895536660167907921591089967922046243014967296;
            6'd20: xpb[28] = 256'd4523128485832663883733241601930416354379124113601674831545181101308436807680;
            6'd21: xpb[28] = 256'd4749284910124297077919903682026937172098080319281758573122440156373858648064;
            6'd22: xpb[28] = 256'd4975441334415930272106565762123457989817036524961842314699699211439280488448;
            6'd23: xpb[28] = 256'd5201597758707563466293227842219978807535992730641926056276958266504702328832;
            6'd24: xpb[28] = 256'd5427754182999196660479889922316499625254948936322009797854217321570124169216;
            6'd25: xpb[28] = 256'd5653910607290829854666552002413020442973905142002093539431476376635546009600;
            6'd26: xpb[28] = 256'd5880067031582463048853214082509541260692861347682177281008735431700967849984;
            6'd27: xpb[28] = 256'd6106223455874096243039876162606062078411817553362261022585994486766389690368;
            6'd28: xpb[28] = 256'd6332379880165729437226538242702582896130773759042344764163253541831811530752;
            6'd29: xpb[28] = 256'd6558536304457362631413200322799103713849729964722428505740512596897233371136;
            6'd30: xpb[28] = 256'd6784692728748995825599862402895624531568686170402512247317771651962655211520;
            6'd31: xpb[28] = 256'd7010849153040629019786524482992145349287642376082595988895030707028077051904;
            6'd32: xpb[28] = 256'd7237005577332262213973186563088666167006598581762679730472289762093498892288;
            6'd33: xpb[28] = 256'd7463162001623895408159848643185186984725554787442763472049548817158920732672;
            6'd34: xpb[28] = 256'd7689318425915528602346510723281707802444510993122847213626807872224342573056;
            6'd35: xpb[28] = 256'd7915474850207161796533172803378228620163467198802930955204066927289764413440;
            6'd36: xpb[28] = 256'd8141631274498794990719834883474749437882423404483014696781325982355186253824;
            6'd37: xpb[28] = 256'd8367787698790428184906496963571270255601379610163098438358585037420608094208;
            6'd38: xpb[28] = 256'd8593944123082061379093159043667791073320335815843182179935844092486029934592;
            6'd39: xpb[28] = 256'd8820100547373694573279821123764311891039292021523265921513103147551451774976;
            6'd40: xpb[28] = 256'd9046256971665327767466483203860832708758248227203349663090362202616873615360;
            6'd41: xpb[28] = 256'd9272413395956960961653145283957353526477204432883433404667621257682295455744;
            6'd42: xpb[28] = 256'd9498569820248594155839807364053874344196160638563517146244880312747717296128;
            6'd43: xpb[28] = 256'd9724726244540227350026469444150395161915116844243600887822139367813139136512;
            6'd44: xpb[28] = 256'd9950882668831860544213131524246915979634073049923684629399398422878560976896;
            6'd45: xpb[28] = 256'd10177039093123493738399793604343436797353029255603768370976657477943982817280;
            6'd46: xpb[28] = 256'd10403195517415126932586455684439957615071985461283852112553916533009404657664;
            6'd47: xpb[28] = 256'd10629351941706760126773117764536478432790941666963935854131175588074826498048;
            6'd48: xpb[28] = 256'd10855508365998393320959779844632999250509897872644019595708434643140248338432;
            6'd49: xpb[28] = 256'd11081664790290026515146441924729520068228854078324103337285693698205670178816;
            6'd50: xpb[28] = 256'd11307821214581659709333104004826040885947810284004187078862952753271092019200;
            6'd51: xpb[28] = 256'd11533977638873292903519766084922561703666766489684270820440211808336513859584;
            6'd52: xpb[28] = 256'd11760134063164926097706428165019082521385722695364354562017470863401935699968;
            6'd53: xpb[28] = 256'd11986290487456559291893090245115603339104678901044438303594729918467357540352;
            6'd54: xpb[28] = 256'd12212446911748192486079752325212124156823635106724522045171988973532779380736;
            6'd55: xpb[28] = 256'd12438603336039825680266414405308644974542591312404605786749248028598201221120;
            6'd56: xpb[28] = 256'd12664759760331458874453076485405165792261547518084689528326507083663623061504;
            6'd57: xpb[28] = 256'd12890916184623092068639738565501686609980503723764773269903766138729044901888;
            6'd58: xpb[28] = 256'd13117072608914725262826400645598207427699459929444857011481025193794466742272;
            6'd59: xpb[28] = 256'd13343229033206358457013062725694728245418416135124940753058284248859888582656;
            6'd60: xpb[28] = 256'd13569385457497991651199724805791249063137372340805024494635543303925310423040;
            6'd61: xpb[28] = 256'd13795541881789624845386386885887769880856328546485108236212802358990732263424;
            6'd62: xpb[28] = 256'd14021698306081258039573048965984290698575284752165191977790061414056154103808;
            6'd63: xpb[28] = 256'd14247854730372891233759711046080811516294240957845275719367320469121575944192;
        endcase
    end

    always_comb begin
        case(flag[29])
            6'd0: xpb[29] = 256'd0;
            6'd1: xpb[29] = 256'd14474011154664524427946373126177332334013197163525359460944579524186997784576;
            6'd2: xpb[29] = 256'd28948022309329048855892746252354664668026394327050718921889159048373995569152;
            6'd3: xpb[29] = 256'd43422033463993573283839119378531997002039591490576078382833738572560993353728;
            6'd4: xpb[29] = 256'd57896044618658097711785492504709329336052788654101437843778318096747991138304;
            6'd5: xpb[29] = 256'd72370055773322622139731865630886661670065985817626797304722897620934988922880;
            6'd6: xpb[29] = 256'd86844066927987146567678238757063994004079182981152156765667477145121986707456;
            6'd7: xpb[29] = 256'd101318078082651670995624611883241326338092380144677516226612056669308984492032;
            6'd8: xpb[29] = 256'd26959946667150639795397765905855223316278684233135442260206297284609;
            6'd9: xpb[29] = 256'd14474011181624471095097012921575098239868420479804043694080021784393295069185;
            6'd10: xpb[29] = 256'd28948022336288995523043386047752430573881617643329403155024601308580292853761;
            6'd11: xpb[29] = 256'd43422033490953519950989759173929762907894814806854762615969180832767290638337;
            6'd12: xpb[29] = 256'd57896044645618044378936132300107095241908011970380122076913760356954288422913;
            6'd13: xpb[29] = 256'd72370055800282568806882505426284427575921209133905481537858339881141286207489;
            6'd14: xpb[29] = 256'd86844066954947093234828878552461759909934406297430840998802919405328283992065;
            6'd15: xpb[29] = 256'd101318078109611617662775251678639092243947603460956200459747498929515281776641;
            6'd16: xpb[29] = 256'd53919893334301279590795531811710446632557368466270884520412594569218;
            6'd17: xpb[29] = 256'd14474011208584417762247652716972864145723643796082727927215464044599592353794;
            6'd18: xpb[29] = 256'd28948022363248942190194025843150196479736840959608087388160043568786590138370;
            6'd19: xpb[29] = 256'd43422033517913466618140398969327528813750038123133446849104623092973587922946;
            6'd20: xpb[29] = 256'd57896044672577991046086772095504861147763235286658806310049202617160585707522;
            6'd21: xpb[29] = 256'd72370055827242515474033145221682193481776432450184165770993782141347583492098;
            6'd22: xpb[29] = 256'd86844066981907039901979518347859525815789629613709525231938361665534581276674;
            6'd23: xpb[29] = 256'd101318078136571564329925891474036858149802826777234884692882941189721579061250;
            6'd24: xpb[29] = 256'd80879840001451919386193297717565669948836052699406326780618891853827;
            6'd25: xpb[29] = 256'd14474011235544364429398292512370630051578867112361412160350906304805889638403;
            6'd26: xpb[29] = 256'd28948022390208888857344665638547962385592064275886771621295485828992887422979;
            6'd27: xpb[29] = 256'd43422033544873413285291038764725294719605261439412131082240065353179885207555;
            6'd28: xpb[29] = 256'd57896044699537937713237411890902627053618458602937490543184644877366882992131;
            6'd29: xpb[29] = 256'd72370055854202462141183785017079959387631655766462850004129224401553880776707;
            6'd30: xpb[29] = 256'd86844067008866986569130158143257291721644852929988209465073803925740878561283;
            6'd31: xpb[29] = 256'd101318078163531510997076531269434624055658050093513568926018383449927876345859;
            6'd32: xpb[29] = 256'd107839786668602559181591063623420893265114736932541769040825189138436;
            6'd33: xpb[29] = 256'd14474011262504311096548932307768395957434090428640096393486348565012186923012;
            6'd34: xpb[29] = 256'd28948022417168835524495305433945728291447287592165455854430928089199184707588;
            6'd35: xpb[29] = 256'd43422033571833359952441678560123060625460484755690815315375507613386182492164;
            6'd36: xpb[29] = 256'd57896044726497884380388051686300392959473681919216174776320087137573180276740;
            6'd37: xpb[29] = 256'd72370055881162408808334424812477725293486879082741534237264666661760178061316;
            6'd38: xpb[29] = 256'd86844067035826933236280797938655057627500076246266893698209246185947175845892;
            6'd39: xpb[29] = 256'd101318078190491457664227171064832389961513273409792253159153825710134173630468;
            6'd40: xpb[29] = 256'd134799733335753198976988829529276116581393421165677211301031486423045;
            6'd41: xpb[29] = 256'd14474011289464257763699572103166161863289313744918780626621790825218484207621;
            6'd42: xpb[29] = 256'd28948022444128782191645945229343494197302510908444140087566370349405481992197;
            6'd43: xpb[29] = 256'd43422033598793306619592318355520826531315708071969499548510949873592479776773;
            6'd44: xpb[29] = 256'd57896044753457831047538691481698158865328905235494859009455529397779477561349;
            6'd45: xpb[29] = 256'd72370055908122355475485064607875491199342102399020218470400108921966475345925;
            6'd46: xpb[29] = 256'd86844067062786879903431437734052823533355299562545577931344688446153473130501;
            6'd47: xpb[29] = 256'd101318078217451404331377810860230155867368496726070937392289267970340470915077;
            6'd48: xpb[29] = 256'd161759680002903838772386595435131339897672105398812653561237783707654;
            6'd49: xpb[29] = 256'd14474011316424204430850211898563927769144537061197464859757233085424781492230;
            6'd50: xpb[29] = 256'd28948022471088728858796585024741260103157734224722824320701812609611779276806;
            6'd51: xpb[29] = 256'd43422033625753253286742958150918592437170931388248183781646392133798777061382;
            6'd52: xpb[29] = 256'd57896044780417777714689331277095924771184128551773543242590971657985774845958;
            6'd53: xpb[29] = 256'd72370055935082302142635704403273257105197325715298902703535551182172772630534;
            6'd54: xpb[29] = 256'd86844067089746826570582077529450589439210522878824262164480130706359770415110;
            6'd55: xpb[29] = 256'd101318078244411350998528450655627921773223720042349621625424710230546768199686;
            6'd56: xpb[29] = 256'd188719626670054478567784361340986563213950789631948095821444080992263;
            6'd57: xpb[29] = 256'd14474011343384151098000851693961693674999760377476149092892675345631078776839;
            6'd58: xpb[29] = 256'd28948022498048675525947224820139026009012957541001508553837254869818076561415;
            6'd59: xpb[29] = 256'd43422033652713199953893597946316358343026154704526868014781834394005074345991;
            6'd60: xpb[29] = 256'd57896044807377724381839971072493690677039351868052227475726413918192072130567;
            6'd61: xpb[29] = 256'd72370055962042248809786344198671023011052549031577586936670993442379069915143;
            6'd62: xpb[29] = 256'd86844067116706773237732717324848355345065746195102946397615572966566067699719;
            6'd63: xpb[29] = 256'd101318078271371297665679090451025687679078943358628305858560152490753065484295;
        endcase
    end

    always_comb begin
        case(flag[30])
            6'd0: xpb[30] = 256'd0;
            6'd1: xpb[30] = 256'd53919893334301279590795531811710446632557368466270884520412594569218;
            6'd2: xpb[30] = 256'd107839786668602559181591063623420893265114736932541769040825189138436;
            6'd3: xpb[30] = 256'd161759680002903838772386595435131339897672105398812653561237783707654;
            6'd4: xpb[30] = 256'd215679573337205118363182127246841786530229473865083538081650378276872;
            6'd5: xpb[30] = 256'd269599466671506397953977659058552233162786842331354422602062972846090;
            6'd6: xpb[30] = 256'd323519360005807677544773190870262679795344210797625307122475567415308;
            6'd7: xpb[30] = 256'd377439253340108957135568722681973126427901579263896191642888161984526;
            6'd8: xpb[30] = 256'd431359146674410236726364254493683573060458947730167076163300756553744;
            6'd9: xpb[30] = 256'd485279040008711516317159786305394019693016316196437960683713351122962;
            6'd10: xpb[30] = 256'd539198933343012795907955318117104466325573684662708845204125945692180;
            6'd11: xpb[30] = 256'd593118826677314075498750849928814912958131053128979729724538540261398;
            6'd12: xpb[30] = 256'd647038720011615355089546381740525359590688421595250614244951134830616;
            6'd13: xpb[30] = 256'd700958613345916634680341913552235806223245790061521498765363729399834;
            6'd14: xpb[30] = 256'd754878506680217914271137445363946252855803158527792383285776323969052;
            6'd15: xpb[30] = 256'd808798400014519193861932977175656699488360526994063267806188918538270;
            6'd16: xpb[30] = 256'd862718293348820473452728508987367146120917895460334152326601513107488;
            6'd17: xpb[30] = 256'd916638186683121753043524040799077592753475263926605036847014107676706;
            6'd18: xpb[30] = 256'd970558080017423032634319572610788039386032632392875921367426702245924;
            6'd19: xpb[30] = 256'd1024477973351724312225115104422498486018590000859146805887839296815142;
            6'd20: xpb[30] = 256'd1078397866686025591815910636234208932651147369325417690408251891384360;
            6'd21: xpb[30] = 256'd1132317760020326871406706168045919379283704737791688574928664485953578;
            6'd22: xpb[30] = 256'd1186237653354628150997501699857629825916262106257959459449077080522796;
            6'd23: xpb[30] = 256'd1240157546688929430588297231669340272548819474724230343969489675092014;
            6'd24: xpb[30] = 256'd1294077440023230710179092763481050719181376843190501228489902269661232;
            6'd25: xpb[30] = 256'd1347997333357531989769888295292761165813934211656772113010314864230450;
            6'd26: xpb[30] = 256'd1401917226691833269360683827104471612446491580123042997530727458799668;
            6'd27: xpb[30] = 256'd1455837120026134548951479358916182059079048948589313882051140053368886;
            6'd28: xpb[30] = 256'd1509757013360435828542274890727892505711606317055584766571552647938104;
            6'd29: xpb[30] = 256'd1563676906694737108133070422539602952344163685521855651091965242507322;
            6'd30: xpb[30] = 256'd1617596800029038387723865954351313398976721053988126535612377837076540;
            6'd31: xpb[30] = 256'd1671516693363339667314661486163023845609278422454397420132790431645758;
            6'd32: xpb[30] = 256'd1725436586697640946905457017974734292241835790920668304653203026214976;
            6'd33: xpb[30] = 256'd1779356480031942226496252549786444738874393159386939189173615620784194;
            6'd34: xpb[30] = 256'd1833276373366243506087048081598155185506950527853210073694028215353412;
            6'd35: xpb[30] = 256'd1887196266700544785677843613409865632139507896319480958214440809922630;
            6'd36: xpb[30] = 256'd1941116160034846065268639145221576078772065264785751842734853404491848;
            6'd37: xpb[30] = 256'd1995036053369147344859434677033286525404622633252022727255265999061066;
            6'd38: xpb[30] = 256'd2048955946703448624450230208844996972037180001718293611775678593630284;
            6'd39: xpb[30] = 256'd2102875840037749904041025740656707418669737370184564496296091188199502;
            6'd40: xpb[30] = 256'd2156795733372051183631821272468417865302294738650835380816503782768720;
            6'd41: xpb[30] = 256'd2210715626706352463222616804280128311934852107117106265336916377337938;
            6'd42: xpb[30] = 256'd2264635520040653742813412336091838758567409475583377149857328971907156;
            6'd43: xpb[30] = 256'd2318555413374955022404207867903549205199966844049648034377741566476374;
            6'd44: xpb[30] = 256'd2372475306709256301995003399715259651832524212515918918898154161045592;
            6'd45: xpb[30] = 256'd2426395200043557581585798931526970098465081580982189803418566755614810;
            6'd46: xpb[30] = 256'd2480315093377858861176594463338680545097638949448460687938979350184028;
            6'd47: xpb[30] = 256'd2534234986712160140767389995150390991730196317914731572459391944753246;
            6'd48: xpb[30] = 256'd2588154880046461420358185526962101438362753686381002456979804539322464;
            6'd49: xpb[30] = 256'd2642074773380762699948981058773811884995311054847273341500217133891682;
            6'd50: xpb[30] = 256'd2695994666715063979539776590585522331627868423313544226020629728460900;
            6'd51: xpb[30] = 256'd2749914560049365259130572122397232778260425791779815110541042323030118;
            6'd52: xpb[30] = 256'd2803834453383666538721367654208943224892983160246085995061454917599336;
            6'd53: xpb[30] = 256'd2857754346717967818312163186020653671525540528712356879581867512168554;
            6'd54: xpb[30] = 256'd2911674240052269097902958717832364118158097897178627764102280106737772;
            6'd55: xpb[30] = 256'd2965594133386570377493754249644074564790655265644898648622692701306990;
            6'd56: xpb[30] = 256'd3019514026720871657084549781455785011423212634111169533143105295876208;
            6'd57: xpb[30] = 256'd3073433920055172936675345313267495458055770002577440417663517890445426;
            6'd58: xpb[30] = 256'd3127353813389474216266140845079205904688327371043711302183930485014644;
            6'd59: xpb[30] = 256'd3181273706723775495856936376890916351320884739509982186704343079583862;
            6'd60: xpb[30] = 256'd3235193600058076775447731908702626797953442107976253071224755674153080;
            6'd61: xpb[30] = 256'd3289113493392378055038527440514337244585999476442523955745168268722298;
            6'd62: xpb[30] = 256'd3343033386726679334629322972326047691218556844908794840265580863291516;
            6'd63: xpb[30] = 256'd3396953280060980614220118504137758137851114213375065724785993457860734;
        endcase
    end

    always_comb begin
        case(flag[31])
            6'd0: xpb[31] = 256'd0;
            6'd1: xpb[31] = 256'd3450873173395281893810914035949468584483671581841336609306406052429952;
            6'd2: xpb[31] = 256'd6901746346790563787621828071898937168967343163682673218612812104859904;
            6'd3: xpb[31] = 256'd10352619520185845681432742107848405753451014745524009827919218157289856;
            6'd4: xpb[31] = 256'd13803492693581127575243656143797874337934686327365346437225624209719808;
            6'd5: xpb[31] = 256'd17254365866976409469054570179747342922418357909206683046532030262149760;
            6'd6: xpb[31] = 256'd20705239040371691362865484215696811506902029491048019655838436314579712;
            6'd7: xpb[31] = 256'd24156112213766973256676398251646280091385701072889356265144842367009664;
            6'd8: xpb[31] = 256'd27606985387162255150487312287595748675869372654730692874451248419439616;
            6'd9: xpb[31] = 256'd31057858560557537044298226323545217260353044236572029483757654471869568;
            6'd10: xpb[31] = 256'd34508731733952818938109140359494685844836715818413366093064060524299520;
            6'd11: xpb[31] = 256'd37959604907348100831920054395444154429320387400254702702370466576729472;
            6'd12: xpb[31] = 256'd41410478080743382725730968431393623013804058982096039311676872629159424;
            6'd13: xpb[31] = 256'd44861351254138664619541882467343091598287730563937375920983278681589376;
            6'd14: xpb[31] = 256'd48312224427533946513352796503292560182771402145778712530289684734019328;
            6'd15: xpb[31] = 256'd51763097600929228407163710539242028767255073727620049139596090786449280;
            6'd16: xpb[31] = 256'd55213970774324510300974624575191497351738745309461385748902496838879232;
            6'd17: xpb[31] = 256'd58664843947719792194785538611140965936222416891302722358208902891309184;
            6'd18: xpb[31] = 256'd62115717121115074088596452647090434520706088473144058967515308943739136;
            6'd19: xpb[31] = 256'd65566590294510355982407366683039903105189760054985395576821714996169088;
            6'd20: xpb[31] = 256'd69017463467905637876218280718989371689673431636826732186128121048599040;
            6'd21: xpb[31] = 256'd72468336641300919770029194754938840274157103218668068795434527101028992;
            6'd22: xpb[31] = 256'd75919209814696201663840108790888308858640774800509405404740933153458944;
            6'd23: xpb[31] = 256'd79370082988091483557651022826837777443124446382350742014047339205888896;
            6'd24: xpb[31] = 256'd82820956161486765451461936862787246027608117964192078623353745258318848;
            6'd25: xpb[31] = 256'd86271829334882047345272850898736714612091789546033415232660151310748800;
            6'd26: xpb[31] = 256'd89722702508277329239083764934686183196575461127874751841966557363178752;
            6'd27: xpb[31] = 256'd93173575681672611132894678970635651781059132709716088451272963415608704;
            6'd28: xpb[31] = 256'd96624448855067893026705593006585120365542804291557425060579369468038656;
            6'd29: xpb[31] = 256'd100075322028463174920516507042534588950026475873398761669885775520468608;
            6'd30: xpb[31] = 256'd103526195201858456814327421078484057534510147455240098279192181572898560;
            6'd31: xpb[31] = 256'd106977068375253738708138335114433526118993819037081434888498587625328512;
            6'd32: xpb[31] = 256'd110427941548649020601949249150382994703477490618922771497804993677758464;
            6'd33: xpb[31] = 256'd113878814722044302495760163186332463287961162200764108107111399730188416;
            6'd34: xpb[31] = 256'd117329687895439584389571077222281931872444833782605444716417805782618368;
            6'd35: xpb[31] = 256'd120780561068834866283381991258231400456928505364446781325724211835048320;
            6'd36: xpb[31] = 256'd124231434242230148177192905294180869041412176946288117935030617887478272;
            6'd37: xpb[31] = 256'd127682307415625430071003819330130337625895848528129454544337023939908224;
            6'd38: xpb[31] = 256'd131133180589020711964814733366079806210379520109970791153643429992338176;
            6'd39: xpb[31] = 256'd134584053762415993858625647402029274794863191691812127762949836044768128;
            6'd40: xpb[31] = 256'd138034926935811275752436561437978743379346863273653464372256242097198080;
            6'd41: xpb[31] = 256'd141485800109206557646247475473928211963830534855494800981562648149628032;
            6'd42: xpb[31] = 256'd144936673282601839540058389509877680548314206437336137590869054202057984;
            6'd43: xpb[31] = 256'd148387546455997121433869303545827149132797878019177474200175460254487936;
            6'd44: xpb[31] = 256'd151838419629392403327680217581776617717281549601018810809481866306917888;
            6'd45: xpb[31] = 256'd155289292802787685221491131617726086301765221182860147418788272359347840;
            6'd46: xpb[31] = 256'd158740165976182967115302045653675554886248892764701484028094678411777792;
            6'd47: xpb[31] = 256'd162191039149578249009112959689625023470732564346542820637401084464207744;
            6'd48: xpb[31] = 256'd165641912322973530902923873725574492055216235928384157246707490516637696;
            6'd49: xpb[31] = 256'd169092785496368812796734787761523960639699907510225493856013896569067648;
            6'd50: xpb[31] = 256'd172543658669764094690545701797473429224183579092066830465320302621497600;
            6'd51: xpb[31] = 256'd175994531843159376584356615833422897808667250673908167074626708673927552;
            6'd52: xpb[31] = 256'd179445405016554658478167529869372366393150922255749503683933114726357504;
            6'd53: xpb[31] = 256'd182896278189949940371978443905321834977634593837590840293239520778787456;
            6'd54: xpb[31] = 256'd186347151363345222265789357941271303562118265419432176902545926831217408;
            6'd55: xpb[31] = 256'd189798024536740504159600271977220772146601937001273513511852332883647360;
            6'd56: xpb[31] = 256'd193248897710135786053411186013170240731085608583114850121158738936077312;
            6'd57: xpb[31] = 256'd196699770883531067947222100049119709315569280164956186730465144988507264;
            6'd58: xpb[31] = 256'd200150644056926349841033014085069177900052951746797523339771551040937216;
            6'd59: xpb[31] = 256'd203601517230321631734843928121018646484536623328638859949077957093367168;
            6'd60: xpb[31] = 256'd207052390403716913628654842156968115069020294910480196558384363145797120;
            6'd61: xpb[31] = 256'd210503263577112195522465756192917583653503966492321533167690769198227072;
            6'd62: xpb[31] = 256'd213954136750507477416276670228867052237987638074162869776997175250657024;
            6'd63: xpb[31] = 256'd217405009923902759310087584264816520822471309656004206386303581303086976;
        endcase
    end

    always_comb begin
        case(flag[32])
            6'd0: xpb[32] = 256'd0;
            6'd1: xpb[32] = 256'd220855883097298041203898498300765989406954981237845542995609987355516928;
            6'd2: xpb[32] = 256'd441711766194596082407796996601531978813909962475691085991219974711033856;
            6'd3: xpb[32] = 256'd662567649291894123611695494902297968220864943713536628986829962066550784;
            6'd4: xpb[32] = 256'd883423532389192164815593993203063957627819924951382171982439949422067712;
            6'd5: xpb[32] = 256'd1104279415486490206019492491503829947034774906189227714978049936777584640;
            6'd6: xpb[32] = 256'd1325135298583788247223390989804595936441729887427073257973659924133101568;
            6'd7: xpb[32] = 256'd1545991181681086288427289488105361925848684868664918800969269911488618496;
            6'd8: xpb[32] = 256'd1766847064778384329631187986406127915255639849902764343964879898844135424;
            6'd9: xpb[32] = 256'd1987702947875682370835086484706893904662594831140609886960489886199652352;
            6'd10: xpb[32] = 256'd2208558830972980412038984983007659894069549812378455429956099873555169280;
            6'd11: xpb[32] = 256'd2429414714070278453242883481308425883476504793616300972951709860910686208;
            6'd12: xpb[32] = 256'd2650270597167576494446781979609191872883459774854146515947319848266203136;
            6'd13: xpb[32] = 256'd2871126480264874535650680477909957862290414756091992058942929835621720064;
            6'd14: xpb[32] = 256'd3091982363362172576854578976210723851697369737329837601938539822977236992;
            6'd15: xpb[32] = 256'd3312838246459470618058477474511489841104324718567683144934149810332753920;
            6'd16: xpb[32] = 256'd3533694129556768659262375972812255830511279699805528687929759797688270848;
            6'd17: xpb[32] = 256'd3754550012654066700466274471113021819918234681043374230925369785043787776;
            6'd18: xpb[32] = 256'd3975405895751364741670172969413787809325189662281219773920979772399304704;
            6'd19: xpb[32] = 256'd4196261778848662782874071467714553798732144643519065316916589759754821632;
            6'd20: xpb[32] = 256'd4417117661945960824077969966015319788139099624756910859912199747110338560;
            6'd21: xpb[32] = 256'd4637973545043258865281868464316085777546054605994756402907809734465855488;
            6'd22: xpb[32] = 256'd4858829428140556906485766962616851766953009587232601945903419721821372416;
            6'd23: xpb[32] = 256'd5079685311237854947689665460917617756359964568470447488899029709176889344;
            6'd24: xpb[32] = 256'd5300541194335152988893563959218383745766919549708293031894639696532406272;
            6'd25: xpb[32] = 256'd5521397077432451030097462457519149735173874530946138574890249683887923200;
            6'd26: xpb[32] = 256'd5742252960529749071301360955819915724580829512183984117885859671243440128;
            6'd27: xpb[32] = 256'd5963108843627047112505259454120681713987784493421829660881469658598957056;
            6'd28: xpb[32] = 256'd6183964726724345153709157952421447703394739474659675203877079645954473984;
            6'd29: xpb[32] = 256'd6404820609821643194913056450722213692801694455897520746872689633309990912;
            6'd30: xpb[32] = 256'd6625676492918941236116954949022979682208649437135366289868299620665507840;
            6'd31: xpb[32] = 256'd6846532376016239277320853447323745671615604418373211832863909608021024768;
            6'd32: xpb[32] = 256'd7067388259113537318524751945624511661022559399611057375859519595376541696;
            6'd33: xpb[32] = 256'd7288244142210835359728650443925277650429514380848902918855129582732058624;
            6'd34: xpb[32] = 256'd7509100025308133400932548942226043639836469362086748461850739570087575552;
            6'd35: xpb[32] = 256'd7729955908405431442136447440526809629243424343324594004846349557443092480;
            6'd36: xpb[32] = 256'd7950811791502729483340345938827575618650379324562439547841959544798609408;
            6'd37: xpb[32] = 256'd8171667674600027524544244437128341608057334305800285090837569532154126336;
            6'd38: xpb[32] = 256'd8392523557697325565748142935429107597464289287038130633833179519509643264;
            6'd39: xpb[32] = 256'd8613379440794623606952041433729873586871244268275976176828789506865160192;
            6'd40: xpb[32] = 256'd8834235323891921648155939932030639576278199249513821719824399494220677120;
            6'd41: xpb[32] = 256'd9055091206989219689359838430331405565685154230751667262820009481576194048;
            6'd42: xpb[32] = 256'd9275947090086517730563736928632171555092109211989512805815619468931710976;
            6'd43: xpb[32] = 256'd9496802973183815771767635426932937544499064193227358348811229456287227904;
            6'd44: xpb[32] = 256'd9717658856281113812971533925233703533906019174465203891806839443642744832;
            6'd45: xpb[32] = 256'd9938514739378411854175432423534469523312974155703049434802449430998261760;
            6'd46: xpb[32] = 256'd10159370622475709895379330921835235512719929136940894977798059418353778688;
            6'd47: xpb[32] = 256'd10380226505573007936583229420136001502126884118178740520793669405709295616;
            6'd48: xpb[32] = 256'd10601082388670305977787127918436767491533839099416586063789279393064812544;
            6'd49: xpb[32] = 256'd10821938271767604018991026416737533480940794080654431606784889380420329472;
            6'd50: xpb[32] = 256'd11042794154864902060194924915038299470347749061892277149780499367775846400;
            6'd51: xpb[32] = 256'd11263650037962200101398823413339065459754704043130122692776109355131363328;
            6'd52: xpb[32] = 256'd11484505921059498142602721911639831449161659024367968235771719342486880256;
            6'd53: xpb[32] = 256'd11705361804156796183806620409940597438568614005605813778767329329842397184;
            6'd54: xpb[32] = 256'd11926217687254094225010518908241363427975568986843659321762939317197914112;
            6'd55: xpb[32] = 256'd12147073570351392266214417406542129417382523968081504864758549304553431040;
            6'd56: xpb[32] = 256'd12367929453448690307418315904842895406789478949319350407754159291908947968;
            6'd57: xpb[32] = 256'd12588785336545988348622214403143661396196433930557195950749769279264464896;
            6'd58: xpb[32] = 256'd12809641219643286389826112901444427385603388911795041493745379266619981824;
            6'd59: xpb[32] = 256'd13030497102740584431030011399745193375010343893032887036740989253975498752;
            6'd60: xpb[32] = 256'd13251352985837882472233909898045959364417298874270732579736599241331015680;
            6'd61: xpb[32] = 256'd13472208868935180513437808396346725353824253855508578122732209228686532608;
            6'd62: xpb[32] = 256'd13693064752032478554641706894647491343231208836746423665727819216042049536;
            6'd63: xpb[32] = 256'd13913920635129776595845605392948257332638163817984269208723429203397566464;
        endcase
    end

    always_comb begin
        case(flag[33])
            6'd0: xpb[33] = 256'd0;
            6'd1: xpb[33] = 256'd3533694129556768659262375972812255830511279699805528687929759797688270848;
            6'd2: xpb[33] = 256'd7067388259113537318524751945624511661022559399611057375859519595376541696;
            6'd3: xpb[33] = 256'd10601082388670305977787127918436767491533839099416586063789279393064812544;
            6'd4: xpb[33] = 256'd14134776518227074637049503891249023322045118799222114751719039190753083392;
            6'd5: xpb[33] = 256'd17668470647783843296311879864061279152556398499027643439648798988441354240;
            6'd6: xpb[33] = 256'd21202164777340611955574255836873534983067678198833172127578558786129625088;
            6'd7: xpb[33] = 256'd24735858906897380614836631809685790813578957898638700815508318583817895936;
            6'd8: xpb[33] = 256'd28269553036454149274099007782498046644090237598444229503438078381506166784;
            6'd9: xpb[33] = 256'd31803247166010917933361383755310302474601517298249758191367838179194437632;
            6'd10: xpb[33] = 256'd35336941295567686592623759728122558305112796998055286879297597976882708480;
            6'd11: xpb[33] = 256'd38870635425124455251886135700934814135624076697860815567227357774570979328;
            6'd12: xpb[33] = 256'd42404329554681223911148511673747069966135356397666344255157117572259250176;
            6'd13: xpb[33] = 256'd45938023684237992570410887646559325796646636097471872943086877369947521024;
            6'd14: xpb[33] = 256'd49471717813794761229673263619371581627157915797277401631016637167635791872;
            6'd15: xpb[33] = 256'd53005411943351529888935639592183837457669195497082930318946396965324062720;
            6'd16: xpb[33] = 256'd56539106072908298548198015564996093288180475196888459006876156763012333568;
            6'd17: xpb[33] = 256'd60072800202465067207460391537808349118691754896693987694805916560700604416;
            6'd18: xpb[33] = 256'd63606494332021835866722767510620604949203034596499516382735676358388875264;
            6'd19: xpb[33] = 256'd67140188461578604525985143483432860779714314296305045070665436156077146112;
            6'd20: xpb[33] = 256'd70673882591135373185247519456245116610225593996110573758595195953765416960;
            6'd21: xpb[33] = 256'd74207576720692141844509895429057372440736873695916102446524955751453687808;
            6'd22: xpb[33] = 256'd77741270850248910503772271401869628271248153395721631134454715549141958656;
            6'd23: xpb[33] = 256'd81274964979805679163034647374681884101759433095527159822384475346830229504;
            6'd24: xpb[33] = 256'd84808659109362447822297023347494139932270712795332688510314235144518500352;
            6'd25: xpb[33] = 256'd88342353238919216481559399320306395762781992495138217198243994942206771200;
            6'd26: xpb[33] = 256'd91876047368475985140821775293118651593293272194943745886173754739895042048;
            6'd27: xpb[33] = 256'd95409741498032753800084151265930907423804551894749274574103514537583312896;
            6'd28: xpb[33] = 256'd98943435627589522459346527238743163254315831594554803262033274335271583744;
            6'd29: xpb[33] = 256'd102477129757146291118608903211555419084827111294360331949963034132959854592;
            6'd30: xpb[33] = 256'd106010823886703059777871279184367674915338390994165860637892793930648125440;
            6'd31: xpb[33] = 256'd109544518016259828437133655157179930745849670693971389325822553728336396288;
            6'd32: xpb[33] = 256'd113078212145816597096396031129992186576360950393776918013752313526024667136;
            6'd33: xpb[33] = 256'd116611906275373365755658407102804442406872230093582446701682073323712937984;
            6'd34: xpb[33] = 256'd120145600404930134414920783075616698237383509793387975389611833121401208832;
            6'd35: xpb[33] = 256'd123679294534486903074183159048428954067894789493193504077541592919089479680;
            6'd36: xpb[33] = 256'd127212988664043671733445535021241209898406069192999032765471352716777750528;
            6'd37: xpb[33] = 256'd130746682793600440392707910994053465728917348892804561453401112514466021376;
            6'd38: xpb[33] = 256'd134280376923157209051970286966865721559428628592610090141330872312154292224;
            6'd39: xpb[33] = 256'd137814071052713977711232662939677977389939908292415618829260632109842563072;
            6'd40: xpb[33] = 256'd141347765182270746370495038912490233220451187992221147517190391907530833920;
            6'd41: xpb[33] = 256'd144881459311827515029757414885302489050962467692026676205120151705219104768;
            6'd42: xpb[33] = 256'd148415153441384283689019790858114744881473747391832204893049911502907375616;
            6'd43: xpb[33] = 256'd151948847570941052348282166830927000711985027091637733580979671300595646464;
            6'd44: xpb[33] = 256'd155482541700497821007544542803739256542496306791443262268909431098283917312;
            6'd45: xpb[33] = 256'd159016235830054589666806918776551512373007586491248790956839190895972188160;
            6'd46: xpb[33] = 256'd162549929959611358326069294749363768203518866191054319644768950693660459008;
            6'd47: xpb[33] = 256'd166083624089168126985331670722176024034030145890859848332698710491348729856;
            6'd48: xpb[33] = 256'd169617318218724895644594046694988279864541425590665377020628470289037000704;
            6'd49: xpb[33] = 256'd173151012348281664303856422667800535695052705290470905708558230086725271552;
            6'd50: xpb[33] = 256'd176684706477838432963118798640612791525563984990276434396487989884413542400;
            6'd51: xpb[33] = 256'd180218400607395201622381174613425047356075264690081963084417749682101813248;
            6'd52: xpb[33] = 256'd183752094736951970281643550586237303186586544389887491772347509479790084096;
            6'd53: xpb[33] = 256'd187285788866508738940905926559049559017097824089693020460277269277478354944;
            6'd54: xpb[33] = 256'd190819482996065507600168302531861814847609103789498549148207029075166625792;
            6'd55: xpb[33] = 256'd194353177125622276259430678504674070678120383489304077836136788872854896640;
            6'd56: xpb[33] = 256'd197886871255179044918693054477486326508631663189109606524066548670543167488;
            6'd57: xpb[33] = 256'd201420565384735813577955430450298582339142942888915135211996308468231438336;
            6'd58: xpb[33] = 256'd204954259514292582237217806423110838169654222588720663899926068265919709184;
            6'd59: xpb[33] = 256'd208487953643849350896480182395923094000165502288526192587855828063607980032;
            6'd60: xpb[33] = 256'd212021647773406119555742558368735349830676781988331721275785587861296250880;
            6'd61: xpb[33] = 256'd215555341902962888215004934341547605661188061688137249963715347658984521728;
            6'd62: xpb[33] = 256'd219089036032519656874267310314359861491699341387942778651645107456672792576;
            6'd63: xpb[33] = 256'd222622730162076425533529686287172117322210621087748307339574867254361063424;
        endcase
    end

    always_comb begin
        case(flag[34])
            6'd0: xpb[34] = 256'd0;
            6'd1: xpb[34] = 256'd226156424291633194192792062259984373152721900787553836027504627052049334272;
            6'd2: xpb[34] = 256'd452312848583266388385584124519968746305443801575107672055009254104098668544;
            6'd3: xpb[34] = 256'd678469272874899582578376186779953119458165702362661508082513881156148002816;
            6'd4: xpb[34] = 256'd904625697166532776771168249039937492610887603150215344110018508208197337088;
            6'd5: xpb[34] = 256'd1130782121458165970963960311299921865763609503937769180137523135260246671360;
            6'd6: xpb[34] = 256'd1356938545749799165156752373559906238916331404725323016165027762312296005632;
            6'd7: xpb[34] = 256'd1583094970041432359349544435819890612069053305512876852192532389364345339904;
            6'd8: xpb[34] = 256'd1809251394333065553542336498079874985221775206300430688220037016416394674176;
            6'd9: xpb[34] = 256'd2035407818624698747735128560339859358374497107087984524247541643468444008448;
            6'd10: xpb[34] = 256'd2261564242916331941927920622599843731527219007875538360275046270520493342720;
            6'd11: xpb[34] = 256'd2487720667207965136120712684859828104679940908663092196302550897572542676992;
            6'd12: xpb[34] = 256'd2713877091499598330313504747119812477832662809450646032330055524624592011264;
            6'd13: xpb[34] = 256'd2940033515791231524506296809379796850985384710238199868357560151676641345536;
            6'd14: xpb[34] = 256'd3166189940082864718699088871639781224138106611025753704385064778728690679808;
            6'd15: xpb[34] = 256'd3392346364374497912891880933899765597290828511813307540412569405780740014080;
            6'd16: xpb[34] = 256'd3618502788666131107084672996159749970443550412600861376440074032832789348352;
            6'd17: xpb[34] = 256'd3844659212957764301277465058419734343596272313388415212467578659884838682624;
            6'd18: xpb[34] = 256'd4070815637249397495470257120679718716748994214175969048495083286936888016896;
            6'd19: xpb[34] = 256'd4296972061541030689663049182939703089901716114963522884522587913988937351168;
            6'd20: xpb[34] = 256'd4523128485832663883855841245199687463054438015751076720550092541040986685440;
            6'd21: xpb[34] = 256'd4749284910124297078048633307459671836207159916538630556577597168093036019712;
            6'd22: xpb[34] = 256'd4975441334415930272241425369719656209359881817326184392605101795145085353984;
            6'd23: xpb[34] = 256'd5201597758707563466434217431979640582512603718113738228632606422197134688256;
            6'd24: xpb[34] = 256'd5427754182999196660627009494239624955665325618901292064660111049249184022528;
            6'd25: xpb[34] = 256'd5653910607290829854819801556499609328818047519688845900687615676301233356800;
            6'd26: xpb[34] = 256'd5880067031582463049012593618759593701970769420476399736715120303353282691072;
            6'd27: xpb[34] = 256'd6106223455874096243205385681019578075123491321263953572742624930405332025344;
            6'd28: xpb[34] = 256'd6332379880165729437398177743279562448276213222051507408770129557457381359616;
            6'd29: xpb[34] = 256'd6558536304457362631590969805539546821428935122839061244797634184509430693888;
            6'd30: xpb[34] = 256'd6784692728748995825783761867799531194581657023626615080825138811561480028160;
            6'd31: xpb[34] = 256'd7010849153040629019976553930059515567734378924414168916852643438613529362432;
            6'd32: xpb[34] = 256'd7237005577332262214169345992319499940887100825201722752880148065665578696704;
            6'd33: xpb[34] = 256'd7463162001623895408362138054579484314039822725989276588907652692717628030976;
            6'd34: xpb[34] = 256'd7689318425915528602554930116839468687192544626776830424935157319769677365248;
            6'd35: xpb[34] = 256'd7915474850207161796747722179099453060345266527564384260962661946821726699520;
            6'd36: xpb[34] = 256'd8141631274498794990940514241359437433497988428351938096990166573873776033792;
            6'd37: xpb[34] = 256'd8367787698790428185133306303619421806650710329139491933017671200925825368064;
            6'd38: xpb[34] = 256'd8593944123082061379326098365879406179803432229927045769045175827977874702336;
            6'd39: xpb[34] = 256'd8820100547373694573518890428139390552956154130714599605072680455029924036608;
            6'd40: xpb[34] = 256'd9046256971665327767711682490399374926108876031502153441100185082081973370880;
            6'd41: xpb[34] = 256'd9272413395956960961904474552659359299261597932289707277127689709134022705152;
            6'd42: xpb[34] = 256'd9498569820248594156097266614919343672414319833077261113155194336186072039424;
            6'd43: xpb[34] = 256'd9724726244540227350290058677179328045567041733864814949182698963238121373696;
            6'd44: xpb[34] = 256'd9950882668831860544482850739439312418719763634652368785210203590290170707968;
            6'd45: xpb[34] = 256'd10177039093123493738675642801699296791872485535439922621237708217342220042240;
            6'd46: xpb[34] = 256'd10403195517415126932868434863959281165025207436227476457265212844394269376512;
            6'd47: xpb[34] = 256'd10629351941706760127061226926219265538177929337015030293292717471446318710784;
            6'd48: xpb[34] = 256'd10855508365998393321254018988479249911330651237802584129320222098498368045056;
            6'd49: xpb[34] = 256'd11081664790290026515446811050739234284483373138590137965347726725550417379328;
            6'd50: xpb[34] = 256'd11307821214581659709639603112999218657636095039377691801375231352602466713600;
            6'd51: xpb[34] = 256'd11533977638873292903832395175259203030788816940165245637402735979654516047872;
            6'd52: xpb[34] = 256'd11760134063164926098025187237519187403941538840952799473430240606706565382144;
            6'd53: xpb[34] = 256'd11986290487456559292217979299779171777094260741740353309457745233758614716416;
            6'd54: xpb[34] = 256'd12212446911748192486410771362039156150246982642527907145485249860810664050688;
            6'd55: xpb[34] = 256'd12438603336039825680603563424299140523399704543315460981512754487862713384960;
            6'd56: xpb[34] = 256'd12664759760331458874796355486559124896552426444103014817540259114914762719232;
            6'd57: xpb[34] = 256'd12890916184623092068989147548819109269705148344890568653567763741966812053504;
            6'd58: xpb[34] = 256'd13117072608914725263181939611079093642857870245678122489595268369018861387776;
            6'd59: xpb[34] = 256'd13343229033206358457374731673339078016010592146465676325622772996070910722048;
            6'd60: xpb[34] = 256'd13569385457497991651567523735599062389163314047253230161650277623122960056320;
            6'd61: xpb[34] = 256'd13795541881789624845760315797859046762316035948040783997677782250175009390592;
            6'd62: xpb[34] = 256'd14021698306081258039953107860119031135468757848828337833705286877227058724864;
            6'd63: xpb[34] = 256'd14247854730372891234145899922379015508621479749615891669732791504279108059136;
        endcase
    end

    always_comb begin
        case(flag[35])
            6'd0: xpb[35] = 256'd0;
            6'd1: xpb[35] = 256'd14474011154664524428338691984638999881774201650403445505760296131331157393408;
            6'd2: xpb[35] = 256'd28948022309329048856677383969277999763548403300806891011520592262662314786816;
            6'd3: xpb[35] = 256'd43422033463993573285016075953916999645322604951210336517280888393993472180224;
            6'd4: xpb[35] = 256'd57896044618658097713354767938555999527096806601613782023041184525324629573632;
            6'd5: xpb[35] = 256'd72370055773322622141693459923194999408871008252017227528801480656655786967040;
            6'd6: xpb[35] = 256'd86844066927987146570032151907833999290645209902420673034561776787986944360448;
            6'd7: xpb[35] = 256'd101318078082651670998370843892472999172419411552824118540322072919318101753856;
            6'd8: xpb[35] = 256'd26959946670289190663091106287943259211303372591661175117359574155265;
            6'd9: xpb[35] = 256'd14474011181624471098627882647730106169717460861706818097421471248690731548673;
            6'd10: xpb[35] = 256'd28948022336288995526966574632369106051491662512110263603181767380021888942081;
            6'd11: xpb[35] = 256'd43422033490953519955305266617008105933265864162513709108942063511353046335489;
            6'd12: xpb[35] = 256'd57896044645618044383643958601647105815040065812917154614702359642684203728897;
            6'd13: xpb[35] = 256'd72370055800282568811982650586286105696814267463320600120462655774015361122305;
            6'd14: xpb[35] = 256'd86844066954947093240321342570925105578588469113724045626222951905346518515713;
            6'd15: xpb[35] = 256'd101318078109611617668660034555564105460362670764127491131983248036677675909121;
            6'd16: xpb[35] = 256'd53919893340578381326182212575886518422606745183322350234719148310530;
            6'd17: xpb[35] = 256'd14474011208584417768917073310821212457660720073010190689082646366050305703938;
            6'd18: xpb[35] = 256'd28948022363248942197255765295460212339434921723413636194842942497381463097346;
            6'd19: xpb[35] = 256'd43422033517913466625594457280099212221209123373817081700603238628712620490754;
            6'd20: xpb[35] = 256'd57896044672577991053933149264738212102983325024220527206363534760043777884162;
            6'd21: xpb[35] = 256'd72370055827242515482271841249377211984757526674623972712123830891374935277570;
            6'd22: xpb[35] = 256'd86844066981907039910610533234016211866531728325027418217884127022706092670978;
            6'd23: xpb[35] = 256'd101318078136571564338949225218655211748305929975430863723644423154037250064386;
            6'd24: xpb[35] = 256'd80879840010867571989273318863829777633910117774983525352078722465795;
            6'd25: xpb[35] = 256'd14474011235544364439206263973912318745603979284313563280743821483409879859203;
            6'd26: xpb[35] = 256'd28948022390208888867544955958551318627378180934717008786504117614741037252611;
            6'd27: xpb[35] = 256'd43422033544873413295883647943190318509152382585120454292264413746072194646019;
            6'd28: xpb[35] = 256'd57896044699537937724222339927829318390926584235523899798024709877403352039427;
            6'd29: xpb[35] = 256'd72370055854202462152561031912468318272700785885927345303785006008734509432835;
            6'd30: xpb[35] = 256'd86844067008866986580899723897107318154474987536330790809545302140065666826243;
            6'd31: xpb[35] = 256'd101318078163531511009238415881746318036249189186734236315305598271396824219651;
            6'd32: xpb[35] = 256'd107839786681156762652364425151773036845213490366644700469438296621060;
            6'd33: xpb[35] = 256'd14474011262504311109495454637003425033547238495616935872404996600769454014468;
            6'd34: xpb[35] = 256'd28948022417168835537834146621642424915321440146020381378165292732100611407876;
            6'd35: xpb[35] = 256'd43422033571833359966172838606281424797095641796423826883925588863431768801284;
            6'd36: xpb[35] = 256'd57896044726497884394511530590920424678869843446827272389685884994762926194692;
            6'd37: xpb[35] = 256'd72370055881162408822850222575559424560644045097230717895446181126094083588100;
            6'd38: xpb[35] = 256'd86844067035826933251188914560198424442418246747634163401206477257425240981508;
            6'd39: xpb[35] = 256'd101318078190491457679527606544837424324192448398037608906966773388756398374916;
            6'd40: xpb[35] = 256'd134799733351445953315455531439716296056516862958305875586797870776325;
            6'd41: xpb[35] = 256'd14474011289464257779784645300094531321490497706920308464066171718129028169733;
            6'd42: xpb[35] = 256'd28948022444128782208123337284733531203264699357323753969826467849460185563141;
            6'd43: xpb[35] = 256'd43422033598793306636462029269372531085038901007727199475586763980791342956549;
            6'd44: xpb[35] = 256'd57896044753457831064800721254011530966813102658130644981347060112122500349957;
            6'd45: xpb[35] = 256'd72370055908122355493139413238650530848587304308534090487107356243453657743365;
            6'd46: xpb[35] = 256'd86844067062786879921478105223289530730361505958937535992867652374784815136773;
            6'd47: xpb[35] = 256'd101318078217451404349816797207928530612135707609340981498627948506115972530181;
            6'd48: xpb[35] = 256'd161759680021735143978546637727659555267820235549967050704157444931590;
            6'd49: xpb[35] = 256'd14474011316424204450073835963185637609433756918223681055727346835488602324998;
            6'd50: xpb[35] = 256'd28948022471088728878412527947824637491207958568627126561487642966819759718406;
            6'd51: xpb[35] = 256'd43422033625753253306751219932463637372982160219030572067247939098150917111814;
            6'd52: xpb[35] = 256'd57896044780417777735089911917102637254756361869434017573008235229482074505222;
            6'd53: xpb[35] = 256'd72370055935082302163428603901741637136530563519837463078768531360813231898630;
            6'd54: xpb[35] = 256'd86844067089746826591767295886380637018304765170240908584528827492144389292038;
            6'd55: xpb[35] = 256'd101318078244411351020105987871019636900078966820644354090289123623475546685446;
            6'd56: xpb[35] = 256'd188719626692024334641637744015602814479123608141628225821517019086855;
            6'd57: xpb[35] = 256'd14474011343384151120363026626276743897377016129527053647388521952848176480263;
            6'd58: xpb[35] = 256'd28948022498048675548701718610915743779151217779930499153148818084179333873671;
            6'd59: xpb[35] = 256'd43422033652713199977040410595554743660925419430333944658909114215510491267079;
            6'd60: xpb[35] = 256'd57896044807377724405379102580193743542699621080737390164669410346841648660487;
            6'd61: xpb[35] = 256'd72370055962042248833717794564832743424473822731140835670429706478172806053895;
            6'd62: xpb[35] = 256'd86844067116706773262056486549471743306248024381544281176190002609503963447303;
            6'd63: xpb[35] = 256'd101318078271371297690395178534110743188022226031947726681950298740835120840711;
        endcase
    end

    always_comb begin
        case(flag[36])
            6'd0: xpb[36] = 256'd0;
            6'd1: xpb[36] = 256'd53919893340578381326182212575886518422606745183322350234719148310530;
            6'd2: xpb[36] = 256'd107839786681156762652364425151773036845213490366644700469438296621060;
            6'd3: xpb[36] = 256'd161759680021735143978546637727659555267820235549967050704157444931590;
            6'd4: xpb[36] = 256'd215679573362313525304728850303546073690426980733289400938876593242120;
            6'd5: xpb[36] = 256'd269599466702891906630911062879432592113033725916611751173595741552650;
            6'd6: xpb[36] = 256'd323519360043470287957093275455319110535640471099934101408314889863180;
            6'd7: xpb[36] = 256'd377439253384048669283275488031205628958247216283256451643034038173710;
            6'd8: xpb[36] = 256'd431359146724627050609457700607092147380853961466578801877753186484240;
            6'd9: xpb[36] = 256'd485279040065205431935639913182978665803460706649901152112472334794770;
            6'd10: xpb[36] = 256'd539198933405783813261822125758865184226067451833223502347191483105300;
            6'd11: xpb[36] = 256'd593118826746362194588004338334751702648674197016545852581910631415830;
            6'd12: xpb[36] = 256'd647038720086940575914186550910638221071280942199868202816629779726360;
            6'd13: xpb[36] = 256'd700958613427518957240368763486524739493887687383190553051348928036890;
            6'd14: xpb[36] = 256'd754878506768097338566550976062411257916494432566512903286068076347420;
            6'd15: xpb[36] = 256'd808798400108675719892733188638297776339101177749835253520787224657950;
            6'd16: xpb[36] = 256'd862718293449254101218915401214184294761707922933157603755506372968480;
            6'd17: xpb[36] = 256'd916638186789832482545097613790070813184314668116479953990225521279010;
            6'd18: xpb[36] = 256'd970558080130410863871279826365957331606921413299802304224944669589540;
            6'd19: xpb[36] = 256'd1024477973470989245197462038941843850029528158483124654459663817900070;
            6'd20: xpb[36] = 256'd1078397866811567626523644251517730368452134903666447004694382966210600;
            6'd21: xpb[36] = 256'd1132317760152146007849826464093616886874741648849769354929102114521130;
            6'd22: xpb[36] = 256'd1186237653492724389176008676669503405297348394033091705163821262831660;
            6'd23: xpb[36] = 256'd1240157546833302770502190889245389923719955139216414055398540411142190;
            6'd24: xpb[36] = 256'd1294077440173881151828373101821276442142561884399736405633259559452720;
            6'd25: xpb[36] = 256'd1347997333514459533154555314397162960565168629583058755867978707763250;
            6'd26: xpb[36] = 256'd1401917226855037914480737526973049478987775374766381106102697856073780;
            6'd27: xpb[36] = 256'd1455837120195616295806919739548935997410382119949703456337417004384310;
            6'd28: xpb[36] = 256'd1509757013536194677133101952124822515832988865133025806572136152694840;
            6'd29: xpb[36] = 256'd1563676906876773058459284164700709034255595610316348156806855301005370;
            6'd30: xpb[36] = 256'd1617596800217351439785466377276595552678202355499670507041574449315900;
            6'd31: xpb[36] = 256'd1671516693557929821111648589852482071100809100682992857276293597626430;
            6'd32: xpb[36] = 256'd1725436586898508202437830802428368589523415845866315207511012745936960;
            6'd33: xpb[36] = 256'd1779356480239086583764013015004255107946022591049637557745731894247490;
            6'd34: xpb[36] = 256'd1833276373579664965090195227580141626368629336232959907980451042558020;
            6'd35: xpb[36] = 256'd1887196266920243346416377440156028144791236081416282258215170190868550;
            6'd36: xpb[36] = 256'd1941116160260821727742559652731914663213842826599604608449889339179080;
            6'd37: xpb[36] = 256'd1995036053601400109068741865307801181636449571782926958684608487489610;
            6'd38: xpb[36] = 256'd2048955946941978490394924077883687700059056316966249308919327635800140;
            6'd39: xpb[36] = 256'd2102875840282556871721106290459574218481663062149571659154046784110670;
            6'd40: xpb[36] = 256'd2156795733623135253047288503035460736904269807332894009388765932421200;
            6'd41: xpb[36] = 256'd2210715626963713634373470715611347255326876552516216359623485080731730;
            6'd42: xpb[36] = 256'd2264635520304292015699652928187233773749483297699538709858204229042260;
            6'd43: xpb[36] = 256'd2318555413644870397025835140763120292172090042882861060092923377352790;
            6'd44: xpb[36] = 256'd2372475306985448778352017353339006810594696788066183410327642525663320;
            6'd45: xpb[36] = 256'd2426395200326027159678199565914893329017303533249505760562361673973850;
            6'd46: xpb[36] = 256'd2480315093666605541004381778490779847439910278432828110797080822284380;
            6'd47: xpb[36] = 256'd2534234987007183922330563991066666365862517023616150461031799970594910;
            6'd48: xpb[36] = 256'd2588154880347762303656746203642552884285123768799472811266519118905440;
            6'd49: xpb[36] = 256'd2642074773688340684982928416218439402707730513982795161501238267215970;
            6'd50: xpb[36] = 256'd2695994667028919066309110628794325921130337259166117511735957415526500;
            6'd51: xpb[36] = 256'd2749914560369497447635292841370212439552944004349439861970676563837030;
            6'd52: xpb[36] = 256'd2803834453710075828961475053946098957975550749532762212205395712147560;
            6'd53: xpb[36] = 256'd2857754347050654210287657266521985476398157494716084562440114860458090;
            6'd54: xpb[36] = 256'd2911674240391232591613839479097871994820764239899406912674834008768620;
            6'd55: xpb[36] = 256'd2965594133731810972940021691673758513243370985082729262909553157079150;
            6'd56: xpb[36] = 256'd3019514027072389354266203904249645031665977730266051613144272305389680;
            6'd57: xpb[36] = 256'd3073433920412967735592386116825531550088584475449373963378991453700210;
            6'd58: xpb[36] = 256'd3127353813753546116918568329401418068511191220632696313613710602010740;
            6'd59: xpb[36] = 256'd3181273707094124498244750541977304586933797965816018663848429750321270;
            6'd60: xpb[36] = 256'd3235193600434702879570932754553191105356404710999341014083148898631800;
            6'd61: xpb[36] = 256'd3289113493775281260897114967129077623779011456182663364317868046942330;
            6'd62: xpb[36] = 256'd3343033387115859642223297179704964142201618201365985714552587195252860;
            6'd63: xpb[36] = 256'd3396953280456438023549479392280850660624224946549308064787306343563390;
        endcase
    end

    always_comb begin
        case(flag[37])
            6'd0: xpb[37] = 256'd0;
            6'd1: xpb[37] = 256'd3450873173797016404875661604856737179046831691732630415022025491873920;
            6'd2: xpb[37] = 256'd6901746347594032809751323209713474358093663383465260830044050983747840;
            6'd3: xpb[37] = 256'd10352619521391049214626984814570211537140495075197891245066076475621760;
            6'd4: xpb[37] = 256'd13803492695188065619502646419426948716187326766930521660088101967495680;
            6'd5: xpb[37] = 256'd17254365868985082024378308024283685895234158458663152075110127459369600;
            6'd6: xpb[37] = 256'd20705239042782098429253969629140423074280990150395782490132152951243520;
            6'd7: xpb[37] = 256'd24156112216579114834129631233997160253327821842128412905154178443117440;
            6'd8: xpb[37] = 256'd27606985390376131239005292838853897432374653533861043320176203934991360;
            6'd9: xpb[37] = 256'd31057858564173147643880954443710634611421485225593673735198229426865280;
            6'd10: xpb[37] = 256'd34508731737970164048756616048567371790468316917326304150220254918739200;
            6'd11: xpb[37] = 256'd37959604911767180453632277653424108969515148609058934565242280410613120;
            6'd12: xpb[37] = 256'd41410478085564196858507939258280846148561980300791564980264305902487040;
            6'd13: xpb[37] = 256'd44861351259361213263383600863137583327608811992524195395286331394360960;
            6'd14: xpb[37] = 256'd48312224433158229668259262467994320506655643684256825810308356886234880;
            6'd15: xpb[37] = 256'd51763097606955246073134924072851057685702475375989456225330382378108800;
            6'd16: xpb[37] = 256'd55213970780752262478010585677707794864749307067722086640352407869982720;
            6'd17: xpb[37] = 256'd58664843954549278882886247282564532043796138759454717055374433361856640;
            6'd18: xpb[37] = 256'd62115717128346295287761908887421269222842970451187347470396458853730560;
            6'd19: xpb[37] = 256'd65566590302143311692637570492278006401889802142919977885418484345604480;
            6'd20: xpb[37] = 256'd69017463475940328097513232097134743580936633834652608300440509837478400;
            6'd21: xpb[37] = 256'd72468336649737344502388893701991480759983465526385238715462535329352320;
            6'd22: xpb[37] = 256'd75919209823534360907264555306848217939030297218117869130484560821226240;
            6'd23: xpb[37] = 256'd79370082997331377312140216911704955118077128909850499545506586313100160;
            6'd24: xpb[37] = 256'd82820956171128393717015878516561692297123960601583129960528611804974080;
            6'd25: xpb[37] = 256'd86271829344925410121891540121418429476170792293315760375550637296848000;
            6'd26: xpb[37] = 256'd89722702518722426526767201726275166655217623985048390790572662788721920;
            6'd27: xpb[37] = 256'd93173575692519442931642863331131903834264455676781021205594688280595840;
            6'd28: xpb[37] = 256'd96624448866316459336518524935988641013311287368513651620616713772469760;
            6'd29: xpb[37] = 256'd100075322040113475741394186540845378192358119060246282035638739264343680;
            6'd30: xpb[37] = 256'd103526195213910492146269848145702115371404950751978912450660764756217600;
            6'd31: xpb[37] = 256'd106977068387707508551145509750558852550451782443711542865682790248091520;
            6'd32: xpb[37] = 256'd110427941561504524956021171355415589729498614135444173280704815739965440;
            6'd33: xpb[37] = 256'd113878814735301541360896832960272326908545445827176803695726841231839360;
            6'd34: xpb[37] = 256'd117329687909098557765772494565129064087592277518909434110748866723713280;
            6'd35: xpb[37] = 256'd120780561082895574170648156169985801266639109210642064525770892215587200;
            6'd36: xpb[37] = 256'd124231434256692590575523817774842538445685940902374694940792917707461120;
            6'd37: xpb[37] = 256'd127682307430489606980399479379699275624732772594107325355814943199335040;
            6'd38: xpb[37] = 256'd131133180604286623385275140984556012803779604285839955770836968691208960;
            6'd39: xpb[37] = 256'd134584053778083639790150802589412749982826435977572586185858994183082880;
            6'd40: xpb[37] = 256'd138034926951880656195026464194269487161873267669305216600881019674956800;
            6'd41: xpb[37] = 256'd141485800125677672599902125799126224340920099361037847015903045166830720;
            6'd42: xpb[37] = 256'd144936673299474689004777787403982961519966931052770477430925070658704640;
            6'd43: xpb[37] = 256'd148387546473271705409653449008839698699013762744503107845947096150578560;
            6'd44: xpb[37] = 256'd151838419647068721814529110613696435878060594436235738260969121642452480;
            6'd45: xpb[37] = 256'd155289292820865738219404772218553173057107426127968368675991147134326400;
            6'd46: xpb[37] = 256'd158740165994662754624280433823409910236154257819700999091013172626200320;
            6'd47: xpb[37] = 256'd162191039168459771029156095428266647415201089511433629506035198118074240;
            6'd48: xpb[37] = 256'd165641912342256787434031757033123384594247921203166259921057223609948160;
            6'd49: xpb[37] = 256'd169092785516053803838907418637980121773294752894898890336079249101822080;
            6'd50: xpb[37] = 256'd172543658689850820243783080242836858952341584586631520751101274593696000;
            6'd51: xpb[37] = 256'd175994531863647836648658741847693596131388416278364151166123300085569920;
            6'd52: xpb[37] = 256'd179445405037444853053534403452550333310435247970096781581145325577443840;
            6'd53: xpb[37] = 256'd182896278211241869458410065057407070489482079661829411996167351069317760;
            6'd54: xpb[37] = 256'd186347151385038885863285726662263807668528911353562042411189376561191680;
            6'd55: xpb[37] = 256'd189798024558835902268161388267120544847575743045294672826211402053065600;
            6'd56: xpb[37] = 256'd193248897732632918673037049871977282026622574737027303241233427544939520;
            6'd57: xpb[37] = 256'd196699770906429935077912711476834019205669406428759933656255453036813440;
            6'd58: xpb[37] = 256'd200150644080226951482788373081690756384716238120492564071277478528687360;
            6'd59: xpb[37] = 256'd203601517254023967887664034686547493563763069812225194486299504020561280;
            6'd60: xpb[37] = 256'd207052390427820984292539696291404230742809901503957824901321529512435200;
            6'd61: xpb[37] = 256'd210503263601618000697415357896260967921856733195690455316343555004309120;
            6'd62: xpb[37] = 256'd213954136775415017102291019501117705100903564887423085731365580496183040;
            6'd63: xpb[37] = 256'd217405009949212033507166681105974442279950396579155716146387605988056960;
        endcase
    end

    always_comb begin
        case(flag[38])
            6'd0: xpb[38] = 256'd0;
            6'd1: xpb[38] = 256'd220855883123009049912042342710831179458997228270888346561409631479930880;
            6'd2: xpb[38] = 256'd441711766246018099824084685421662358917994456541776693122819262959861760;
            6'd3: xpb[38] = 256'd662567649369027149736127028132493538376991684812665039684228894439792640;
            6'd4: xpb[38] = 256'd883423532492036199648169370843324717835988913083553386245638525919723520;
            6'd5: xpb[38] = 256'd1104279415615045249560211713554155897294986141354441732807048157399654400;
            6'd6: xpb[38] = 256'd1325135298738054299472254056264987076753983369625330079368457788879585280;
            6'd7: xpb[38] = 256'd1545991181861063349384296398975818256212980597896218425929867420359516160;
            6'd8: xpb[38] = 256'd1766847064984072399296338741686649435671977826167106772491277051839447040;
            6'd9: xpb[38] = 256'd1987702948107081449208381084397480615130975054437995119052686683319377920;
            6'd10: xpb[38] = 256'd2208558831230090499120423427108311794589972282708883465614096314799308800;
            6'd11: xpb[38] = 256'd2429414714353099549032465769819142974048969510979771812175505946279239680;
            6'd12: xpb[38] = 256'd2650270597476108598944508112529974153507966739250660158736915577759170560;
            6'd13: xpb[38] = 256'd2871126480599117648856550455240805332966963967521548505298325209239101440;
            6'd14: xpb[38] = 256'd3091982363722126698768592797951636512425961195792436851859734840719032320;
            6'd15: xpb[38] = 256'd3312838246845135748680635140662467691884958424063325198421144472198963200;
            6'd16: xpb[38] = 256'd3533694129968144798592677483373298871343955652334213544982554103678894080;
            6'd17: xpb[38] = 256'd3754550013091153848504719826084130050802952880605101891543963735158824960;
            6'd18: xpb[38] = 256'd3975405896214162898416762168794961230261950108875990238105373366638755840;
            6'd19: xpb[38] = 256'd4196261779337171948328804511505792409720947337146878584666782998118686720;
            6'd20: xpb[38] = 256'd4417117662460180998240846854216623589179944565417766931228192629598617600;
            6'd21: xpb[38] = 256'd4637973545583190048152889196927454768638941793688655277789602261078548480;
            6'd22: xpb[38] = 256'd4858829428706199098064931539638285948097939021959543624351011892558479360;
            6'd23: xpb[38] = 256'd5079685311829208147976973882349117127556936250230431970912421524038410240;
            6'd24: xpb[38] = 256'd5300541194952217197889016225059948307015933478501320317473831155518341120;
            6'd25: xpb[38] = 256'd5521397078075226247801058567770779486474930706772208664035240786998272000;
            6'd26: xpb[38] = 256'd5742252961198235297713100910481610665933927935043097010596650418478202880;
            6'd27: xpb[38] = 256'd5963108844321244347625143253192441845392925163313985357158060049958133760;
            6'd28: xpb[38] = 256'd6183964727444253397537185595903273024851922391584873703719469681438064640;
            6'd29: xpb[38] = 256'd6404820610567262447449227938614104204310919619855762050280879312917995520;
            6'd30: xpb[38] = 256'd6625676493690271497361270281324935383769916848126650396842288944397926400;
            6'd31: xpb[38] = 256'd6846532376813280547273312624035766563228914076397538743403698575877857280;
            6'd32: xpb[38] = 256'd7067388259936289597185354966746597742687911304668427089965108207357788160;
            6'd33: xpb[38] = 256'd7288244143059298647097397309457428922146908532939315436526517838837719040;
            6'd34: xpb[38] = 256'd7509100026182307697009439652168260101605905761210203783087927470317649920;
            6'd35: xpb[38] = 256'd7729955909305316746921481994879091281064902989481092129649337101797580800;
            6'd36: xpb[38] = 256'd7950811792428325796833524337589922460523900217751980476210746733277511680;
            6'd37: xpb[38] = 256'd8171667675551334846745566680300753639982897446022868822772156364757442560;
            6'd38: xpb[38] = 256'd8392523558674343896657609023011584819441894674293757169333565996237373440;
            6'd39: xpb[38] = 256'd8613379441797352946569651365722415998900891902564645515894975627717304320;
            6'd40: xpb[38] = 256'd8834235324920361996481693708433247178359889130835533862456385259197235200;
            6'd41: xpb[38] = 256'd9055091208043371046393736051144078357818886359106422209017794890677166080;
            6'd42: xpb[38] = 256'd9275947091166380096305778393854909537277883587377310555579204522157096960;
            6'd43: xpb[38] = 256'd9496802974289389146217820736565740716736880815648198902140614153637027840;
            6'd44: xpb[38] = 256'd9717658857412398196129863079276571896195878043919087248702023785116958720;
            6'd45: xpb[38] = 256'd9938514740535407246041905421987403075654875272189975595263433416596889600;
            6'd46: xpb[38] = 256'd10159370623658416295953947764698234255113872500460863941824843048076820480;
            6'd47: xpb[38] = 256'd10380226506781425345865990107409065434572869728731752288386252679556751360;
            6'd48: xpb[38] = 256'd10601082389904434395778032450119896614031866957002640634947662311036682240;
            6'd49: xpb[38] = 256'd10821938273027443445690074792830727793490864185273528981509071942516613120;
            6'd50: xpb[38] = 256'd11042794156150452495602117135541558972949861413544417328070481573996544000;
            6'd51: xpb[38] = 256'd11263650039273461545514159478252390152408858641815305674631891205476474880;
            6'd52: xpb[38] = 256'd11484505922396470595426201820963221331867855870086194021193300836956405760;
            6'd53: xpb[38] = 256'd11705361805519479645338244163674052511326853098357082367754710468436336640;
            6'd54: xpb[38] = 256'd11926217688642488695250286506384883690785850326627970714316120099916267520;
            6'd55: xpb[38] = 256'd12147073571765497745162328849095714870244847554898859060877529731396198400;
            6'd56: xpb[38] = 256'd12367929454888506795074371191806546049703844783169747407438939362876129280;
            6'd57: xpb[38] = 256'd12588785338011515844986413534517377229162842011440635754000348994356060160;
            6'd58: xpb[38] = 256'd12809641221134524894898455877228208408621839239711524100561758625835991040;
            6'd59: xpb[38] = 256'd13030497104257533944810498219939039588080836467982412447123168257315921920;
            6'd60: xpb[38] = 256'd13251352987380542994722540562649870767539833696253300793684577888795852800;
            6'd61: xpb[38] = 256'd13472208870503552044634582905360701946998830924524189140245987520275783680;
            6'd62: xpb[38] = 256'd13693064753626561094546625248071533126457828152795077486807397151755714560;
            6'd63: xpb[38] = 256'd13913920636749570144458667590782364305916825381065965833368806783235645440;
        endcase
    end

    always_comb begin
        case(flag[39])
            6'd0: xpb[39] = 256'd0;
            6'd1: xpb[39] = 256'd3533694129968144798592677483373298871343955652334213544982554103678894080;
            6'd2: xpb[39] = 256'd7067388259936289597185354966746597742687911304668427089965108207357788160;
            6'd3: xpb[39] = 256'd10601082389904434395778032450119896614031866957002640634947662311036682240;
            6'd4: xpb[39] = 256'd14134776519872579194370709933493195485375822609336854179930216414715576320;
            6'd5: xpb[39] = 256'd17668470649840723992963387416866494356719778261671067724912770518394470400;
            6'd6: xpb[39] = 256'd21202164779808868791556064900239793228063733914005281269895324622073364480;
            6'd7: xpb[39] = 256'd24735858909777013590148742383613092099407689566339494814877878725752258560;
            6'd8: xpb[39] = 256'd28269553039745158388741419866986390970751645218673708359860432829431152640;
            6'd9: xpb[39] = 256'd31803247169713303187334097350359689842095600871007921904842986933110046720;
            6'd10: xpb[39] = 256'd35336941299681447985926774833732988713439556523342135449825541036788940800;
            6'd11: xpb[39] = 256'd38870635429649592784519452317106287584783512175676348994808095140467834880;
            6'd12: xpb[39] = 256'd42404329559617737583112129800479586456127467828010562539790649244146728960;
            6'd13: xpb[39] = 256'd45938023689585882381704807283852885327471423480344776084773203347825623040;
            6'd14: xpb[39] = 256'd49471717819554027180297484767226184198815379132678989629755757451504517120;
            6'd15: xpb[39] = 256'd53005411949522171978890162250599483070159334785013203174738311555183411200;
            6'd16: xpb[39] = 256'd56539106079490316777482839733972781941503290437347416719720865658862305280;
            6'd17: xpb[39] = 256'd60072800209458461576075517217346080812847246089681630264703419762541199360;
            6'd18: xpb[39] = 256'd63606494339426606374668194700719379684191201742015843809685973866220093440;
            6'd19: xpb[39] = 256'd67140188469394751173260872184092678555535157394350057354668527969898987520;
            6'd20: xpb[39] = 256'd70673882599362895971853549667465977426879113046684270899651082073577881600;
            6'd21: xpb[39] = 256'd74207576729331040770446227150839276298223068699018484444633636177256775680;
            6'd22: xpb[39] = 256'd77741270859299185569038904634212575169567024351352697989616190280935669760;
            6'd23: xpb[39] = 256'd81274964989267330367631582117585874040910980003686911534598744384614563840;
            6'd24: xpb[39] = 256'd84808659119235475166224259600959172912254935656021125079581298488293457920;
            6'd25: xpb[39] = 256'd88342353249203619964816937084332471783598891308355338624563852591972352000;
            6'd26: xpb[39] = 256'd91876047379171764763409614567705770654942846960689552169546406695651246080;
            6'd27: xpb[39] = 256'd95409741509139909562002292051079069526286802613023765714528960799330140160;
            6'd28: xpb[39] = 256'd98943435639108054360594969534452368397630758265357979259511514903009034240;
            6'd29: xpb[39] = 256'd102477129769076199159187647017825667268974713917692192804494069006687928320;
            6'd30: xpb[39] = 256'd106010823899044343957780324501198966140318669570026406349476623110366822400;
            6'd31: xpb[39] = 256'd109544518029012488756373001984572265011662625222360619894459177214045716480;
            6'd32: xpb[39] = 256'd113078212158980633554965679467945563883006580874694833439441731317724610560;
            6'd33: xpb[39] = 256'd116611906288948778353558356951318862754350536527029046984424285421403504640;
            6'd34: xpb[39] = 256'd120145600418916923152151034434692161625694492179363260529406839525082398720;
            6'd35: xpb[39] = 256'd123679294548885067950743711918065460497038447831697474074389393628761292800;
            6'd36: xpb[39] = 256'd127212988678853212749336389401438759368382403484031687619371947732440186880;
            6'd37: xpb[39] = 256'd130746682808821357547929066884812058239726359136365901164354501836119080960;
            6'd38: xpb[39] = 256'd134280376938789502346521744368185357111070314788700114709337055939797975040;
            6'd39: xpb[39] = 256'd137814071068757647145114421851558655982414270441034328254319610043476869120;
            6'd40: xpb[39] = 256'd141347765198725791943707099334931954853758226093368541799302164147155763200;
            6'd41: xpb[39] = 256'd144881459328693936742299776818305253725102181745702755344284718250834657280;
            6'd42: xpb[39] = 256'd148415153458662081540892454301678552596446137398036968889267272354513551360;
            6'd43: xpb[39] = 256'd151948847588630226339485131785051851467790093050371182434249826458192445440;
            6'd44: xpb[39] = 256'd155482541718598371138077809268425150339134048702705395979232380561871339520;
            6'd45: xpb[39] = 256'd159016235848566515936670486751798449210478004355039609524214934665550233600;
            6'd46: xpb[39] = 256'd162549929978534660735263164235171748081821960007373823069197488769229127680;
            6'd47: xpb[39] = 256'd166083624108502805533855841718545046953165915659708036614180042872908021760;
            6'd48: xpb[39] = 256'd169617318238470950332448519201918345824509871312042250159162596976586915840;
            6'd49: xpb[39] = 256'd173151012368439095131041196685291644695853826964376463704145151080265809920;
            6'd50: xpb[39] = 256'd176684706498407239929633874168664943567197782616710677249127705183944704000;
            6'd51: xpb[39] = 256'd180218400628375384728226551652038242438541738269044890794110259287623598080;
            6'd52: xpb[39] = 256'd183752094758343529526819229135411541309885693921379104339092813391302492160;
            6'd53: xpb[39] = 256'd187285788888311674325411906618784840181229649573713317884075367494981386240;
            6'd54: xpb[39] = 256'd190819483018279819124004584102158139052573605226047531429057921598660280320;
            6'd55: xpb[39] = 256'd194353177148247963922597261585531437923917560878381744974040475702339174400;
            6'd56: xpb[39] = 256'd197886871278216108721189939068904736795261516530715958519023029806018068480;
            6'd57: xpb[39] = 256'd201420565408184253519782616552278035666605472183050172064005583909696962560;
            6'd58: xpb[39] = 256'd204954259538152398318375294035651334537949427835384385608988138013375856640;
            6'd59: xpb[39] = 256'd208487953668120543116967971519024633409293383487718599153970692117054750720;
            6'd60: xpb[39] = 256'd212021647798088687915560649002397932280637339140052812698953246220733644800;
            6'd61: xpb[39] = 256'd215555341928056832714153326485771231151981294792387026243935800324412538880;
            6'd62: xpb[39] = 256'd219089036058024977512746003969144530023325250444721239788918354428091432960;
            6'd63: xpb[39] = 256'd222622730187993122311338681452517828894669206097055453333900908531770327040;
        endcase
    end

    always_comb begin
        case(flag[40])
            6'd0: xpb[40] = 256'd0;
            6'd1: xpb[40] = 256'd226156424317961267109931358935891127766013161749389666878883462635449221120;
            6'd2: xpb[40] = 256'd452312848635922534219862717871782255532026323498779333757766925270898442240;
            6'd3: xpb[40] = 256'd678469272953883801329794076807673383298039485248169000636650387906347663360;
            6'd4: xpb[40] = 256'd904625697271845068439725435743564511064052646997558667515533850541796884480;
            6'd5: xpb[40] = 256'd1130782121589806335549656794679455638830065808746948334394417313177246105600;
            6'd6: xpb[40] = 256'd1356938545907767602659588153615346766596078970496338001273300775812695326720;
            6'd7: xpb[40] = 256'd1583094970225728869769519512551237894362092132245727668152184238448144547840;
            6'd8: xpb[40] = 256'd1809251394543690136879450871487129022128105293995117335031067701083593768960;
            6'd9: xpb[40] = 256'd2035407818861651403989382230423020149894118455744507001909951163719042990080;
            6'd10: xpb[40] = 256'd2261564243179612671099313589358911277660131617493896668788834626354492211200;
            6'd11: xpb[40] = 256'd2487720667497573938209244948294802405426144779243286335667718088989941432320;
            6'd12: xpb[40] = 256'd2713877091815535205319176307230693533192157940992676002546601551625390653440;
            6'd13: xpb[40] = 256'd2940033516133496472429107666166584660958171102742065669425485014260839874560;
            6'd14: xpb[40] = 256'd3166189940451457739539039025102475788724184264491455336304368476896289095680;
            6'd15: xpb[40] = 256'd3392346364769419006648970384038366916490197426240845003183251939531738316800;
            6'd16: xpb[40] = 256'd3618502789087380273758901742974258044256210587990234670062135402167187537920;
            6'd17: xpb[40] = 256'd3844659213405341540868833101910149172022223749739624336941018864802636759040;
            6'd18: xpb[40] = 256'd4070815637723302807978764460846040299788236911489014003819902327438085980160;
            6'd19: xpb[40] = 256'd4296972062041264075088695819781931427554250073238403670698785790073535201280;
            6'd20: xpb[40] = 256'd4523128486359225342198627178717822555320263234987793337577669252708984422400;
            6'd21: xpb[40] = 256'd4749284910677186609308558537653713683086276396737183004456552715344433643520;
            6'd22: xpb[40] = 256'd4975441334995147876418489896589604810852289558486572671335436177979882864640;
            6'd23: xpb[40] = 256'd5201597759313109143528421255525495938618302720235962338214319640615332085760;
            6'd24: xpb[40] = 256'd5427754183631070410638352614461387066384315881985352005093203103250781306880;
            6'd25: xpb[40] = 256'd5653910607949031677748283973397278194150329043734741671972086565886230528000;
            6'd26: xpb[40] = 256'd5880067032266992944858215332333169321916342205484131338850970028521679749120;
            6'd27: xpb[40] = 256'd6106223456584954211968146691269060449682355367233521005729853491157128970240;
            6'd28: xpb[40] = 256'd6332379880902915479078078050204951577448368528982910672608736953792578191360;
            6'd29: xpb[40] = 256'd6558536305220876746188009409140842705214381690732300339487620416428027412480;
            6'd30: xpb[40] = 256'd6784692729538838013297940768076733832980394852481690006366503879063476633600;
            6'd31: xpb[40] = 256'd7010849153856799280407872127012624960746408014231079673245387341698925854720;
            6'd32: xpb[40] = 256'd7237005578174760547517803485948516088512421175980469340124270804334375075840;
            6'd33: xpb[40] = 256'd7463162002492721814627734844884407216278434337729859007003154266969824296960;
            6'd34: xpb[40] = 256'd7689318426810683081737666203820298344044447499479248673882037729605273518080;
            6'd35: xpb[40] = 256'd7915474851128644348847597562756189471810460661228638340760921192240722739200;
            6'd36: xpb[40] = 256'd8141631275446605615957528921692080599576473822978028007639804654876171960320;
            6'd37: xpb[40] = 256'd8367787699764566883067460280627971727342486984727417674518688117511621181440;
            6'd38: xpb[40] = 256'd8593944124082528150177391639563862855108500146476807341397571580147070402560;
            6'd39: xpb[40] = 256'd8820100548400489417287322998499753982874513308226197008276455042782519623680;
            6'd40: xpb[40] = 256'd9046256972718450684397254357435645110640526469975586675155338505417968844800;
            6'd41: xpb[40] = 256'd9272413397036411951507185716371536238406539631724976342034221968053418065920;
            6'd42: xpb[40] = 256'd9498569821354373218617117075307427366172552793474366008913105430688867287040;
            6'd43: xpb[40] = 256'd9724726245672334485727048434243318493938565955223755675791988893324316508160;
            6'd44: xpb[40] = 256'd9950882669990295752836979793179209621704579116973145342670872355959765729280;
            6'd45: xpb[40] = 256'd10177039094308257019946911152115100749470592278722535009549755818595214950400;
            6'd46: xpb[40] = 256'd10403195518626218287056842511050991877236605440471924676428639281230664171520;
            6'd47: xpb[40] = 256'd10629351942944179554166773869986883005002618602221314343307522743866113392640;
            6'd48: xpb[40] = 256'd10855508367262140821276705228922774132768631763970704010186406206501562613760;
            6'd49: xpb[40] = 256'd11081664791580102088386636587858665260534644925720093677065289669137011834880;
            6'd50: xpb[40] = 256'd11307821215898063355496567946794556388300658087469483343944173131772461056000;
            6'd51: xpb[40] = 256'd11533977640216024622606499305730447516066671249218873010823056594407910277120;
            6'd52: xpb[40] = 256'd11760134064533985889716430664666338643832684410968262677701940057043359498240;
            6'd53: xpb[40] = 256'd11986290488851947156826362023602229771598697572717652344580823519678808719360;
            6'd54: xpb[40] = 256'd12212446913169908423936293382538120899364710734467042011459706982314257940480;
            6'd55: xpb[40] = 256'd12438603337487869691046224741474012027130723896216431678338590444949707161600;
            6'd56: xpb[40] = 256'd12664759761805830958156156100409903154896737057965821345217473907585156382720;
            6'd57: xpb[40] = 256'd12890916186123792225266087459345794282662750219715211012096357370220605603840;
            6'd58: xpb[40] = 256'd13117072610441753492376018818281685410428763381464600678975240832856054824960;
            6'd59: xpb[40] = 256'd13343229034759714759485950177217576538194776543213990345854124295491504046080;
            6'd60: xpb[40] = 256'd13569385459077676026595881536153467665960789704963380012733007758126953267200;
            6'd61: xpb[40] = 256'd13795541883395637293705812895089358793726802866712769679611891220762402488320;
            6'd62: xpb[40] = 256'd14021698307713598560815744254025249921492816028462159346490774683397851709440;
            6'd63: xpb[40] = 256'd14247854732031559827925675612961141049258829190211549013369658146033300930560;
        endcase
    end

    always_comb begin
        case(flag[41])
            6'd0: xpb[41] = 256'd0;
            6'd1: xpb[41] = 256'd14474011156349521095035606971897032177024842351960938680248541608668750151680;
            6'd2: xpb[41] = 256'd28948022312699042190071213943794064354049684703921877360497083217337500303360;
            6'd3: xpb[41] = 256'd43422033469048563285106820915691096531074527055882816040745624826006250455040;
            6'd4: xpb[41] = 256'd57896044625398084380142427887588128708099369407843754720994166434675000606720;
            6'd5: xpb[41] = 256'd72370055781747605475178034859485160885124211759804693401242708043343750758400;
            6'd6: xpb[41] = 256'd86844066938097126570213641831382193062149054111765632081491249652012500910080;
            6'd7: xpb[41] = 256'd101318078094446647665249248803279225239173896463726570761739791260681251061760;
            6'd8: xpb[41] = 256'd40439920003864510561155364649948384823763317987567138936060316221441;
            6'd9: xpb[41] = 256'd14474011196789441098900117533052396826973227175724256667815680544729066373121;
            6'd10: xpb[41] = 256'd28948022353138962193935724504949429003998069527685195348064222153397816524801;
            6'd11: xpb[41] = 256'd43422033509488483288971331476846461181022911879646134028312763762066566676481;
            6'd12: xpb[41] = 256'd57896044665838004384006938448743493358047754231607072708561305370735316828161;
            6'd13: xpb[41] = 256'd72370055822187525479042545420640525535072596583568011388809846979404066979841;
            6'd14: xpb[41] = 256'd86844066978537046574078152392537557712097438935528950069058388588072817131521;
            6'd15: xpb[41] = 256'd101318078134886567669113759364434589889122281287489888749306930196741567283201;
            6'd16: xpb[41] = 256'd80879840007729021122310729299896769647526635975134277872120632442882;
            6'd17: xpb[41] = 256'd14474011237229361102764628094207761476921611999487574655382819480789382594562;
            6'd18: xpb[41] = 256'd28948022393578882197800235066104793653946454351448513335631361089458132746242;
            6'd19: xpb[41] = 256'd43422033549928403292835842038001825830971296703409452015879902698126882897922;
            6'd20: xpb[41] = 256'd57896044706277924387871449009898858007996139055370390696128444306795633049602;
            6'd21: xpb[41] = 256'd72370055862627445482907055981795890185020981407331329376376985915464383201282;
            6'd22: xpb[41] = 256'd86844067018976966577942662953692922362045823759292268056625527524133133352962;
            6'd23: xpb[41] = 256'd101318078175326487672978269925589954539070666111253206736874069132801883504642;
            6'd24: xpb[41] = 256'd121319760011593531683466093949845154471289953962701416808180948664323;
            6'd25: xpb[41] = 256'd14474011277669281106629138655363126126869996823250892642949958416849698816003;
            6'd26: xpb[41] = 256'd28948022434018802201664745627260158303894839175211831323198500025518448967683;
            6'd27: xpb[41] = 256'd43422033590368323296700352599157190480919681527172770003447041634187199119363;
            6'd28: xpb[41] = 256'd57896044746717844391735959571054222657944523879133708683695583242855949271043;
            6'd29: xpb[41] = 256'd72370055903067365486771566542951254834969366231094647363944124851524699422723;
            6'd30: xpb[41] = 256'd86844067059416886581807173514848287011994208583055586044192666460193449574403;
            6'd31: xpb[41] = 256'd101318078215766407676842780486745319189019050935016524724441208068862199726083;
            6'd32: xpb[41] = 256'd161759680015458042244621458599793539295053271950268555744241264885764;
            6'd33: xpb[41] = 256'd14474011318109201110493649216518490776818381647014210630517097352910015037444;
            6'd34: xpb[41] = 256'd28948022474458722205529256188415522953843223998975149310765638961578765189124;
            6'd35: xpb[41] = 256'd43422033630808243300564863160312555130868066350936087991014180570247515340804;
            6'd36: xpb[41] = 256'd57896044787157764395600470132209587307892908702897026671262722178916265492484;
            6'd37: xpb[41] = 256'd72370055943507285490636077104106619484917751054857965351511263787585015644164;
            6'd38: xpb[41] = 256'd86844067099856806585671684076003651661942593406818904031759805396253765795844;
            6'd39: xpb[41] = 256'd101318078256206327680707291047900683838967435758779842712008347004922515947524;
            6'd40: xpb[41] = 256'd202199600019322552805776823249741924118816589937835694680301581107205;
            6'd41: xpb[41] = 256'd14474011358549121114358159777673855426766766470777528618084236288970331258885;
            6'd42: xpb[41] = 256'd28948022514898642209393766749570887603791608822738467298332777897639081410565;
            6'd43: xpb[41] = 256'd43422033671248163304429373721467919780816451174699405978581319506307831562245;
            6'd44: xpb[41] = 256'd57896044827597684399464980693364951957841293526660344658829861114976581713925;
            6'd45: xpb[41] = 256'd72370055983947205494500587665261984134866135878621283339078402723645331865605;
            6'd46: xpb[41] = 256'd86844067140296726589536194637159016311890978230582222019326944332314082017285;
            6'd47: xpb[41] = 256'd101318078296646247684571801609056048488915820582543160699575485940982832168965;
            6'd48: xpb[41] = 256'd242639520023187063366932187899690308942579907925402833616361897328646;
            6'd49: xpb[41] = 256'd14474011398989041118222670338829220076715151294540846605651375225030647480326;
            6'd50: xpb[41] = 256'd28948022555338562213258277310726252253739993646501785285899916833699397632006;
            6'd51: xpb[41] = 256'd43422033711688083308293884282623284430764835998462723966148458442368147783686;
            6'd52: xpb[41] = 256'd57896044868037604403329491254520316607789678350423662646397000051036897935366;
            6'd53: xpb[41] = 256'd72370056024387125498365098226417348784814520702384601326645541659705648087046;
            6'd54: xpb[41] = 256'd86844067180736646593400705198314380961839363054345540006894083268374398238726;
            6'd55: xpb[41] = 256'd101318078337086167688436312170211413138864205406306478687142624877043148390406;
            6'd56: xpb[41] = 256'd283079440027051573928087552549638693766343225912969972552422213550087;
            6'd57: xpb[41] = 256'd14474011439428961122087180899984584726663536118304164593218514161090963701767;
            6'd58: xpb[41] = 256'd28948022595778482217122787871881616903688378470265103273467055769759713853447;
            6'd59: xpb[41] = 256'd43422033752128003312158394843778649080713220822226041953715597378428464005127;
            6'd60: xpb[41] = 256'd57896044908477524407194001815675681257738063174186980633964138987097214156807;
            6'd61: xpb[41] = 256'd72370056064827045502229608787572713434762905526147919314212680595765964308487;
            6'd62: xpb[41] = 256'd86844067221176566597265215759469745611787747878108857994461222204434714460167;
            6'd63: xpb[41] = 256'd101318078377526087692300822731366777788812590230069796674709763813103464611847;
        endcase
    end

    always_comb begin
        case(flag[42])
            6'd0: xpb[42] = 256'd0;
            6'd1: xpb[42] = 256'd80879840007729021122310729299896769647526635975134277872120632442882;
            6'd2: xpb[42] = 256'd161759680015458042244621458599793539295053271950268555744241264885764;
            6'd3: xpb[42] = 256'd242639520023187063366932187899690308942579907925402833616361897328646;
            6'd4: xpb[42] = 256'd323519360030916084489242917199587078590106543900537111488482529771528;
            6'd5: xpb[42] = 256'd404399200038645105611553646499483848237633179875671389360603162214410;
            6'd6: xpb[42] = 256'd485279040046374126733864375799380617885159815850805667232723794657292;
            6'd7: xpb[42] = 256'd566158880054103147856175105099277387532686451825939945104844427100174;
            6'd8: xpb[42] = 256'd647038720061832168978485834399174157180213087801074222976965059543056;
            6'd9: xpb[42] = 256'd727918560069561190100796563699070926827739723776208500849085691985938;
            6'd10: xpb[42] = 256'd808798400077290211223107292998967696475266359751342778721206324428820;
            6'd11: xpb[42] = 256'd889678240085019232345418022298864466122792995726477056593326956871702;
            6'd12: xpb[42] = 256'd970558080092748253467728751598761235770319631701611334465447589314584;
            6'd13: xpb[42] = 256'd1051437920100477274590039480898658005417846267676745612337568221757466;
            6'd14: xpb[42] = 256'd1132317760108206295712350210198554775065372903651879890209688854200348;
            6'd15: xpb[42] = 256'd1213197600115935316834660939498451544712899539627014168081809486643230;
            6'd16: xpb[42] = 256'd1294077440123664337956971668798348314360426175602148445953930119086112;
            6'd17: xpb[42] = 256'd1374957280131393359079282398098245084007952811577282723826050751528994;
            6'd18: xpb[42] = 256'd1455837120139122380201593127398141853655479447552417001698171383971876;
            6'd19: xpb[42] = 256'd1536716960146851401323903856698038623303006083527551279570292016414758;
            6'd20: xpb[42] = 256'd1617596800154580422446214585997935392950532719502685557442412648857640;
            6'd21: xpb[42] = 256'd1698476640162309443568525315297832162598059355477819835314533281300522;
            6'd22: xpb[42] = 256'd1779356480170038464690836044597728932245585991452954113186653913743404;
            6'd23: xpb[42] = 256'd1860236320177767485813146773897625701893112627428088391058774546186286;
            6'd24: xpb[42] = 256'd1941116160185496506935457503197522471540639263403222668930895178629168;
            6'd25: xpb[42] = 256'd2021996000193225528057768232497419241188165899378356946803015811072050;
            6'd26: xpb[42] = 256'd2102875840200954549180078961797316010835692535353491224675136443514932;
            6'd27: xpb[42] = 256'd2183755680208683570302389691097212780483219171328625502547257075957814;
            6'd28: xpb[42] = 256'd2264635520216412591424700420397109550130745807303759780419377708400696;
            6'd29: xpb[42] = 256'd2345515360224141612547011149697006319778272443278894058291498340843578;
            6'd30: xpb[42] = 256'd2426395200231870633669321878996903089425799079254028336163618973286460;
            6'd31: xpb[42] = 256'd2507275040239599654791632608296799859073325715229162614035739605729342;
            6'd32: xpb[42] = 256'd2588154880247328675913943337596696628720852351204296891907860238172224;
            6'd33: xpb[42] = 256'd2669034720255057697036254066896593398368378987179431169779980870615106;
            6'd34: xpb[42] = 256'd2749914560262786718158564796196490168015905623154565447652101503057988;
            6'd35: xpb[42] = 256'd2830794400270515739280875525496386937663432259129699725524222135500870;
            6'd36: xpb[42] = 256'd2911674240278244760403186254796283707310958895104834003396342767943752;
            6'd37: xpb[42] = 256'd2992554080285973781525496984096180476958485531079968281268463400386634;
            6'd38: xpb[42] = 256'd3073433920293702802647807713396077246606012167055102559140584032829516;
            6'd39: xpb[42] = 256'd3154313760301431823770118442695974016253538803030236837012704665272398;
            6'd40: xpb[42] = 256'd3235193600309160844892429171995870785901065439005371114884825297715280;
            6'd41: xpb[42] = 256'd3316073440316889866014739901295767555548592074980505392756945930158162;
            6'd42: xpb[42] = 256'd3396953280324618887137050630595664325196118710955639670629066562601044;
            6'd43: xpb[42] = 256'd3477833120332347908259361359895561094843645346930773948501187195043926;
            6'd44: xpb[42] = 256'd3558712960340076929381672089195457864491171982905908226373307827486808;
            6'd45: xpb[42] = 256'd3639592800347805950503982818495354634138698618881042504245428459929690;
            6'd46: xpb[42] = 256'd3720472640355534971626293547795251403786225254856176782117549092372572;
            6'd47: xpb[42] = 256'd3801352480363263992748604277095148173433751890831311059989669724815454;
            6'd48: xpb[42] = 256'd3882232320370993013870915006395044943081278526806445337861790357258336;
            6'd49: xpb[42] = 256'd3963112160378722034993225735694941712728805162781579615733910989701218;
            6'd50: xpb[42] = 256'd4043992000386451056115536464994838482376331798756713893606031622144100;
            6'd51: xpb[42] = 256'd4124871840394180077237847194294735252023858434731848171478152254586982;
            6'd52: xpb[42] = 256'd4205751680401909098360157923594632021671385070706982449350272887029864;
            6'd53: xpb[42] = 256'd4286631520409638119482468652894528791318911706682116727222393519472746;
            6'd54: xpb[42] = 256'd4367511360417367140604779382194425560966438342657251005094514151915628;
            6'd55: xpb[42] = 256'd4448391200425096161727090111494322330613964978632385282966634784358510;
            6'd56: xpb[42] = 256'd4529271040432825182849400840794219100261491614607519560838755416801392;
            6'd57: xpb[42] = 256'd4610150880440554203971711570094115869909018250582653838710876049244274;
            6'd58: xpb[42] = 256'd4691030720448283225094022299394012639556544886557788116582996681687156;
            6'd59: xpb[42] = 256'd4771910560456012246216333028693909409204071522532922394455117314130038;
            6'd60: xpb[42] = 256'd4852790400463741267338643757993806178851598158508056672327237946572920;
            6'd61: xpb[42] = 256'd4933670240471470288460954487293702948499124794483190950199358579015802;
            6'd62: xpb[42] = 256'd5014550080479199309583265216593599718146651430458325228071479211458684;
            6'd63: xpb[42] = 256'd5095429920486928330705575945893496487794178066433459505943599843901566;
        endcase
    end

    always_comb begin
        case(flag[43])
            6'd0: xpb[43] = 256'd0;
            6'd1: xpb[43] = 256'd5176309760494657351827886675193393257441704702408593783815720476344448;
            6'd2: xpb[43] = 256'd10352619520989314703655773350386786514883409404817187567631440952688896;
            6'd3: xpb[43] = 256'd15528929281483972055483660025580179772325114107225781351447161429033344;
            6'd4: xpb[43] = 256'd20705239041978629407311546700773573029766818809634375135262881905377792;
            6'd5: xpb[43] = 256'd25881548802473286759139433375966966287208523512042968919078602381722240;
            6'd6: xpb[43] = 256'd31057858562967944110967320051160359544650228214451562702894322858066688;
            6'd7: xpb[43] = 256'd36234168323462601462795206726353752802091932916860156486710043334411136;
            6'd8: xpb[43] = 256'd41410478083957258814623093401547146059533637619268750270525763810755584;
            6'd9: xpb[43] = 256'd46586787844451916166450980076740539316975342321677344054341484287100032;
            6'd10: xpb[43] = 256'd51763097604946573518278866751933932574417047024085937838157204763444480;
            6'd11: xpb[43] = 256'd56939407365441230870106753427127325831858751726494531621972925239788928;
            6'd12: xpb[43] = 256'd62115717125935888221934640102320719089300456428903125405788645716133376;
            6'd13: xpb[43] = 256'd67292026886430545573762526777514112346742161131311719189604366192477824;
            6'd14: xpb[43] = 256'd72468336646925202925590413452707505604183865833720312973420086668822272;
            6'd15: xpb[43] = 256'd77644646407419860277418300127900898861625570536128906757235807145166720;
            6'd16: xpb[43] = 256'd82820956167914517629246186803094292119067275238537500541051527621511168;
            6'd17: xpb[43] = 256'd87997265928409174981074073478287685376508979940946094324867248097855616;
            6'd18: xpb[43] = 256'd93173575688903832332901960153481078633950684643354688108682968574200064;
            6'd19: xpb[43] = 256'd98349885449398489684729846828674471891392389345763281892498689050544512;
            6'd20: xpb[43] = 256'd103526195209893147036557733503867865148834094048171875676314409526888960;
            6'd21: xpb[43] = 256'd108702504970387804388385620179061258406275798750580469460130130003233408;
            6'd22: xpb[43] = 256'd113878814730882461740213506854254651663717503452989063243945850479577856;
            6'd23: xpb[43] = 256'd119055124491377119092041393529448044921159208155397657027761570955922304;
            6'd24: xpb[43] = 256'd124231434251871776443869280204641438178600912857806250811577291432266752;
            6'd25: xpb[43] = 256'd129407744012366433795697166879834831436042617560214844595393011908611200;
            6'd26: xpb[43] = 256'd134584053772861091147525053555028224693484322262623438379208732384955648;
            6'd27: xpb[43] = 256'd139760363533355748499352940230221617950926026965032032163024452861300096;
            6'd28: xpb[43] = 256'd144936673293850405851180826905415011208367731667440625946840173337644544;
            6'd29: xpb[43] = 256'd150112983054345063203008713580608404465809436369849219730655893813988992;
            6'd30: xpb[43] = 256'd155289292814839720554836600255801797723251141072257813514471614290333440;
            6'd31: xpb[43] = 256'd160465602575334377906664486930995190980692845774666407298287334766677888;
            6'd32: xpb[43] = 256'd165641912335829035258492373606188584238134550477075001082103055243022336;
            6'd33: xpb[43] = 256'd170818222096323692610320260281381977495576255179483594865918775719366784;
            6'd34: xpb[43] = 256'd175994531856818349962148146956575370753017959881892188649734496195711232;
            6'd35: xpb[43] = 256'd181170841617313007313976033631768764010459664584300782433550216672055680;
            6'd36: xpb[43] = 256'd186347151377807664665803920306962157267901369286709376217365937148400128;
            6'd37: xpb[43] = 256'd191523461138302322017631806982155550525343073989117970001181657624744576;
            6'd38: xpb[43] = 256'd196699770898796979369459693657348943782784778691526563784997378101089024;
            6'd39: xpb[43] = 256'd201876080659291636721287580332542337040226483393935157568813098577433472;
            6'd40: xpb[43] = 256'd207052390419786294073115467007735730297668188096343751352628819053777920;
            6'd41: xpb[43] = 256'd212228700180280951424943353682929123555109892798752345136444539530122368;
            6'd42: xpb[43] = 256'd217405009940775608776771240358122516812551597501160938920260260006466816;
            6'd43: xpb[43] = 256'd222581319701270266128599127033315910069993302203569532704075980482811264;
            6'd44: xpb[43] = 256'd227757629461764923480427013708509303327435006905978126487891700959155712;
            6'd45: xpb[43] = 256'd232933939222259580832254900383702696584876711608386720271707421435500160;
            6'd46: xpb[43] = 256'd238110248982754238184082787058896089842318416310795314055523141911844608;
            6'd47: xpb[43] = 256'd243286558743248895535910673734089483099760121013203907839338862388189056;
            6'd48: xpb[43] = 256'd248462868503743552887738560409282876357201825715612501623154582864533504;
            6'd49: xpb[43] = 256'd253639178264238210239566447084476269614643530418021095406970303340877952;
            6'd50: xpb[43] = 256'd258815488024732867591394333759669662872085235120429689190786023817222400;
            6'd51: xpb[43] = 256'd263991797785227524943222220434863056129526939822838282974601744293566848;
            6'd52: xpb[43] = 256'd269168107545722182295050107110056449386968644525246876758417464769911296;
            6'd53: xpb[43] = 256'd274344417306216839646877993785249842644410349227655470542233185246255744;
            6'd54: xpb[43] = 256'd279520727066711496998705880460443235901852053930064064326048905722600192;
            6'd55: xpb[43] = 256'd284697036827206154350533767135636629159293758632472658109864626198944640;
            6'd56: xpb[43] = 256'd289873346587700811702361653810830022416735463334881251893680346675289088;
            6'd57: xpb[43] = 256'd295049656348195469054189540486023415674177168037289845677496067151633536;
            6'd58: xpb[43] = 256'd300225966108690126406017427161216808931618872739698439461311787627977984;
            6'd59: xpb[43] = 256'd305402275869184783757845313836410202189060577442107033245127508104322432;
            6'd60: xpb[43] = 256'd310578585629679441109673200511603595446502282144515627028943228580666880;
            6'd61: xpb[43] = 256'd315754895390174098461501087186796988703943986846924220812758949057011328;
            6'd62: xpb[43] = 256'd320931205150668755813328973861990381961385691549332814596574669533355776;
            6'd63: xpb[43] = 256'd326107514911163413165156860537183775218827396251741408380390390009700224;
        endcase
    end

    always_comb begin
        case(flag[44])
            6'd0: xpb[44] = 256'd0;
            6'd1: xpb[44] = 256'd331283824671658070516984747212377168476269100954150002164206110486044672;
            6'd2: xpb[44] = 256'd662567649343316141033969494424754336952538201908300004328412220972089344;
            6'd3: xpb[44] = 256'd993851474014974211550954241637131505428807302862450006492618331458134016;
            6'd4: xpb[44] = 256'd1325135298686632282067938988849508673905076403816600008656824441944178688;
            6'd5: xpb[44] = 256'd1656419123358290352584923736061885842381345504770750010821030552430223360;
            6'd6: xpb[44] = 256'd1987702948029948423101908483274263010857614605724900012985236662916268032;
            6'd7: xpb[44] = 256'd2318986772701606493618893230486640179333883706679050015149442773402312704;
            6'd8: xpb[44] = 256'd2650270597373264564135877977699017347810152807633200017313648883888357376;
            6'd9: xpb[44] = 256'd2981554422044922634652862724911394516286421908587350019477854994374402048;
            6'd10: xpb[44] = 256'd3312838246716580705169847472123771684762691009541500021642061104860446720;
            6'd11: xpb[44] = 256'd3644122071388238775686832219336148853238960110495650023806267215346491392;
            6'd12: xpb[44] = 256'd3975405896059896846203816966548526021715229211449800025970473325832536064;
            6'd13: xpb[44] = 256'd4306689720731554916720801713760903190191498312403950028134679436318580736;
            6'd14: xpb[44] = 256'd4637973545403212987237786460973280358667767413358100030298885546804625408;
            6'd15: xpb[44] = 256'd4969257370074871057754771208185657527144036514312250032463091657290670080;
            6'd16: xpb[44] = 256'd5300541194746529128271755955398034695620305615266400034627297767776714752;
            6'd17: xpb[44] = 256'd5631825019418187198788740702610411864096574716220550036791503878262759424;
            6'd18: xpb[44] = 256'd5963108844089845269305725449822789032572843817174700038955709988748804096;
            6'd19: xpb[44] = 256'd6294392668761503339822710197035166201049112918128850041119916099234848768;
            6'd20: xpb[44] = 256'd6625676493433161410339694944247543369525382019083000043284122209720893440;
            6'd21: xpb[44] = 256'd6956960318104819480856679691459920538001651120037150045448328320206938112;
            6'd22: xpb[44] = 256'd7288244142776477551373664438672297706477920220991300047612534430692982784;
            6'd23: xpb[44] = 256'd7619527967448135621890649185884674874954189321945450049776740541179027456;
            6'd24: xpb[44] = 256'd7950811792119793692407633933097052043430458422899600051940946651665072128;
            6'd25: xpb[44] = 256'd8282095616791451762924618680309429211906727523853750054105152762151116800;
            6'd26: xpb[44] = 256'd8613379441463109833441603427521806380382996624807900056269358872637161472;
            6'd27: xpb[44] = 256'd8944663266134767903958588174734183548859265725762050058433564983123206144;
            6'd28: xpb[44] = 256'd9275947090806425974475572921946560717335534826716200060597771093609250816;
            6'd29: xpb[44] = 256'd9607230915478084044992557669158937885811803927670350062761977204095295488;
            6'd30: xpb[44] = 256'd9938514740149742115509542416371315054288073028624500064926183314581340160;
            6'd31: xpb[44] = 256'd10269798564821400186026527163583692222764342129578650067090389425067384832;
            6'd32: xpb[44] = 256'd10601082389493058256543511910796069391240611230532800069254595535553429504;
            6'd33: xpb[44] = 256'd10932366214164716327060496658008446559716880331486950071418801646039474176;
            6'd34: xpb[44] = 256'd11263650038836374397577481405220823728193149432441100073583007756525518848;
            6'd35: xpb[44] = 256'd11594933863508032468094466152433200896669418533395250075747213867011563520;
            6'd36: xpb[44] = 256'd11926217688179690538611450899645578065145687634349400077911419977497608192;
            6'd37: xpb[44] = 256'd12257501512851348609128435646857955233621956735303550080075626087983652864;
            6'd38: xpb[44] = 256'd12588785337523006679645420394070332402098225836257700082239832198469697536;
            6'd39: xpb[44] = 256'd12920069162194664750162405141282709570574494937211850084404038308955742208;
            6'd40: xpb[44] = 256'd13251352986866322820679389888495086739050764038166000086568244419441786880;
            6'd41: xpb[44] = 256'd13582636811537980891196374635707463907527033139120150088732450529927831552;
            6'd42: xpb[44] = 256'd13913920636209638961713359382919841076003302240074300090896656640413876224;
            6'd43: xpb[44] = 256'd14245204460881297032230344130132218244479571341028450093060862750899920896;
            6'd44: xpb[44] = 256'd14576488285552955102747328877344595412955840441982600095225068861385965568;
            6'd45: xpb[44] = 256'd14907772110224613173264313624556972581432109542936750097389274971872010240;
            6'd46: xpb[44] = 256'd15239055934896271243781298371769349749908378643890900099553481082358054912;
            6'd47: xpb[44] = 256'd15570339759567929314298283118981726918384647744845050101717687192844099584;
            6'd48: xpb[44] = 256'd15901623584239587384815267866194104086860916845799200103881893303330144256;
            6'd49: xpb[44] = 256'd16232907408911245455332252613406481255337185946753350106046099413816188928;
            6'd50: xpb[44] = 256'd16564191233582903525849237360618858423813455047707500108210305524302233600;
            6'd51: xpb[44] = 256'd16895475058254561596366222107831235592289724148661650110374511634788278272;
            6'd52: xpb[44] = 256'd17226758882926219666883206855043612760765993249615800112538717745274322944;
            6'd53: xpb[44] = 256'd17558042707597877737400191602255989929242262350569950114702923855760367616;
            6'd54: xpb[44] = 256'd17889326532269535807917176349468367097718531451524100116867129966246412288;
            6'd55: xpb[44] = 256'd18220610356941193878434161096680744266194800552478250119031336076732456960;
            6'd56: xpb[44] = 256'd18551894181612851948951145843893121434671069653432400121195542187218501632;
            6'd57: xpb[44] = 256'd18883178006284510019468130591105498603147338754386550123359748297704546304;
            6'd58: xpb[44] = 256'd19214461830956168089985115338317875771623607855340700125523954408190590976;
            6'd59: xpb[44] = 256'd19545745655627826160502100085530252940099876956294850127688160518676635648;
            6'd60: xpb[44] = 256'd19877029480299484231019084832742630108576146057249000129852366629162680320;
            6'd61: xpb[44] = 256'd20208313304971142301536069579955007277052415158203150132016572739648724992;
            6'd62: xpb[44] = 256'd20539597129642800372053054327167384445528684259157300134180778850134769664;
            6'd63: xpb[44] = 256'd20870880954314458442570039074379761614004953360111450136344984960620814336;
        endcase
    end

    always_comb begin
        case(flag[45])
            6'd0: xpb[45] = 256'd0;
            6'd1: xpb[45] = 256'd5300541194746529128271755955398034695620305615266400034627297767776714752;
            6'd2: xpb[45] = 256'd10601082389493058256543511910796069391240611230532800069254595535553429504;
            6'd3: xpb[45] = 256'd15901623584239587384815267866194104086860916845799200103881893303330144256;
            6'd4: xpb[45] = 256'd21202164778986116513087023821592138782481222461065600138509191071106859008;
            6'd5: xpb[45] = 256'd26502705973732645641358779776990173478101528076332000173136488838883573760;
            6'd6: xpb[45] = 256'd31803247168479174769630535732388208173721833691598400207763786606660288512;
            6'd7: xpb[45] = 256'd37103788363225703897902291687786242869342139306864800242391084374437003264;
            6'd8: xpb[45] = 256'd42404329557972233026174047643184277564962444922131200277018382142213718016;
            6'd9: xpb[45] = 256'd47704870752718762154445803598582312260582750537397600311645679909990432768;
            6'd10: xpb[45] = 256'd53005411947465291282717559553980346956203056152664000346272977677767147520;
            6'd11: xpb[45] = 256'd58305953142211820410989315509378381651823361767930400380900275445543862272;
            6'd12: xpb[45] = 256'd63606494336958349539261071464776416347443667383196800415527573213320577024;
            6'd13: xpb[45] = 256'd68907035531704878667532827420174451043063972998463200450154870981097291776;
            6'd14: xpb[45] = 256'd74207576726451407795804583375572485738684278613729600484782168748874006528;
            6'd15: xpb[45] = 256'd79508117921197936924076339330970520434304584228996000519409466516650721280;
            6'd16: xpb[45] = 256'd84808659115944466052348095286368555129924889844262400554036764284427436032;
            6'd17: xpb[45] = 256'd90109200310690995180619851241766589825545195459528800588664062052204150784;
            6'd18: xpb[45] = 256'd95409741505437524308891607197164624521165501074795200623291359819980865536;
            6'd19: xpb[45] = 256'd100710282700184053437163363152562659216785806690061600657918657587757580288;
            6'd20: xpb[45] = 256'd106010823894930582565435119107960693912406112305328000692545955355534295040;
            6'd21: xpb[45] = 256'd111311365089677111693706875063358728608026417920594400727173253123311009792;
            6'd22: xpb[45] = 256'd116611906284423640821978631018756763303646723535860800761800550891087724544;
            6'd23: xpb[45] = 256'd121912447479170169950250386974154797999267029151127200796427848658864439296;
            6'd24: xpb[45] = 256'd127212988673916699078522142929552832694887334766393600831055146426641154048;
            6'd25: xpb[45] = 256'd132513529868663228206793898884950867390507640381660000865682444194417868800;
            6'd26: xpb[45] = 256'd137814071063409757335065654840348902086127945996926400900309741962194583552;
            6'd27: xpb[45] = 256'd143114612258156286463337410795746936781748251612192800934937039729971298304;
            6'd28: xpb[45] = 256'd148415153452902815591609166751144971477368557227459200969564337497748013056;
            6'd29: xpb[45] = 256'd153715694647649344719880922706543006172988862842725601004191635265524727808;
            6'd30: xpb[45] = 256'd159016235842395873848152678661941040868609168457992001038818933033301442560;
            6'd31: xpb[45] = 256'd164316777037142402976424434617339075564229474073258401073446230801078157312;
            6'd32: xpb[45] = 256'd169617318231888932104696190572737110259849779688524801108073528568854872064;
            6'd33: xpb[45] = 256'd174917859426635461232967946528135144955470085303791201142700826336631586816;
            6'd34: xpb[45] = 256'd180218400621381990361239702483533179651090390919057601177328124104408301568;
            6'd35: xpb[45] = 256'd185518941816128519489511458438931214346710696534324001211955421872185016320;
            6'd36: xpb[45] = 256'd190819483010875048617783214394329249042331002149590401246582719639961731072;
            6'd37: xpb[45] = 256'd196120024205621577746054970349727283737951307764856801281210017407738445824;
            6'd38: xpb[45] = 256'd201420565400368106874326726305125318433571613380123201315837315175515160576;
            6'd39: xpb[45] = 256'd206721106595114636002598482260523353129191918995389601350464612943291875328;
            6'd40: xpb[45] = 256'd212021647789861165130870238215921387824812224610656001385091910711068590080;
            6'd41: xpb[45] = 256'd217322188984607694259141994171319422520432530225922401419719208478845304832;
            6'd42: xpb[45] = 256'd222622730179354223387413750126717457216052835841188801454346506246622019584;
            6'd43: xpb[45] = 256'd227923271374100752515685506082115491911673141456455201488973804014398734336;
            6'd44: xpb[45] = 256'd233223812568847281643957262037513526607293447071721601523601101782175449088;
            6'd45: xpb[45] = 256'd238524353763593810772229017992911561302913752686988001558228399549952163840;
            6'd46: xpb[45] = 256'd243824894958340339900500773948309595998534058302254401592855697317728878592;
            6'd47: xpb[45] = 256'd249125436153086869028772529903707630694154363917520801627482995085505593344;
            6'd48: xpb[45] = 256'd254425977347833398157044285859105665389774669532787201662110292853282308096;
            6'd49: xpb[45] = 256'd259726518542579927285316041814503700085394975148053601696737590621059022848;
            6'd50: xpb[45] = 256'd265027059737326456413587797769901734781015280763320001731364888388835737600;
            6'd51: xpb[45] = 256'd270327600932072985541859553725299769476635586378586401765992186156612452352;
            6'd52: xpb[45] = 256'd275628142126819514670131309680697804172255891993852801800619483924389167104;
            6'd53: xpb[45] = 256'd280928683321566043798403065636095838867876197609119201835246781692165881856;
            6'd54: xpb[45] = 256'd286229224516312572926674821591493873563496503224385601869874079459942596608;
            6'd55: xpb[45] = 256'd291529765711059102054946577546891908259116808839652001904501377227719311360;
            6'd56: xpb[45] = 256'd296830306905805631183218333502289942954737114454918401939128674995496026112;
            6'd57: xpb[45] = 256'd302130848100552160311490089457687977650357420070184801973755972763272740864;
            6'd58: xpb[45] = 256'd307431389295298689439761845413086012345977725685451202008383270531049455616;
            6'd59: xpb[45] = 256'd312731930490045218568033601368484047041598031300717602043010568298826170368;
            6'd60: xpb[45] = 256'd318032471684791747696305357323882081737218336915984002077637866066602885120;
            6'd61: xpb[45] = 256'd323333012879538276824577113279280116432838642531250402112265163834379599872;
            6'd62: xpb[45] = 256'd328633554074284805952848869234678151128458948146516802146892461602156314624;
            6'd63: xpb[45] = 256'd333934095269031335081120625190076185824079253761783202181519759369933029376;
        endcase
    end

    always_comb begin
        case(flag[46])
            6'd0: xpb[46] = 256'd0;
            6'd1: xpb[46] = 256'd339234636463777864209392381145474220519699559377049602216147057137709744128;
            6'd2: xpb[46] = 256'd678469272927555728418784762290948441039399118754099204432294114275419488256;
            6'd3: xpb[46] = 256'd1017703909391333592628177143436422661559098678131148806648441171413129232384;
            6'd4: xpb[46] = 256'd1356938545855111456837569524581896882078798237508198408864588228550838976512;
            6'd5: xpb[46] = 256'd1696173182318889321046961905727371102598497796885248011080735285688548720640;
            6'd6: xpb[46] = 256'd2035407818782667185256354286872845323118197356262297613296882342826258464768;
            6'd7: xpb[46] = 256'd2374642455246445049465746668018319543637896915639347215513029399963968208896;
            6'd8: xpb[46] = 256'd2713877091710222913675139049163793764157596475016396817729176457101677953024;
            6'd9: xpb[46] = 256'd3053111728174000777884531430309267984677296034393446419945323514239387697152;
            6'd10: xpb[46] = 256'd3392346364637778642093923811454742205196995593770496022161470571377097441280;
            6'd11: xpb[46] = 256'd3731581001101556506303316192600216425716695153147545624377617628514807185408;
            6'd12: xpb[46] = 256'd4070815637565334370512708573745690646236394712524595226593764685652516929536;
            6'd13: xpb[46] = 256'd4410050274029112234722100954891164866756094271901644828809911742790226673664;
            6'd14: xpb[46] = 256'd4749284910492890098931493336036639087275793831278694431026058799927936417792;
            6'd15: xpb[46] = 256'd5088519546956667963140885717182113307795493390655744033242205857065646161920;
            6'd16: xpb[46] = 256'd5427754183420445827350278098327587528315192950032793635458352914203355906048;
            6'd17: xpb[46] = 256'd5766988819884223691559670479473061748834892509409843237674499971341065650176;
            6'd18: xpb[46] = 256'd6106223456348001555769062860618535969354592068786892839890647028478775394304;
            6'd19: xpb[46] = 256'd6445458092811779419978455241764010189874291628163942442106794085616485138432;
            6'd20: xpb[46] = 256'd6784692729275557284187847622909484410393991187540992044322941142754194882560;
            6'd21: xpb[46] = 256'd7123927365739335148397240004054958630913690746918041646539088199891904626688;
            6'd22: xpb[46] = 256'd7463162002203113012606632385200432851433390306295091248755235257029614370816;
            6'd23: xpb[46] = 256'd7802396638666890876816024766345907071953089865672140850971382314167324114944;
            6'd24: xpb[46] = 256'd8141631275130668741025417147491381292472789425049190453187529371305033859072;
            6'd25: xpb[46] = 256'd8480865911594446605234809528636855512992488984426240055403676428442743603200;
            6'd26: xpb[46] = 256'd8820100548058224469444201909782329733512188543803289657619823485580453347328;
            6'd27: xpb[46] = 256'd9159335184522002333653594290927803954031888103180339259835970542718163091456;
            6'd28: xpb[46] = 256'd9498569820985780197862986672073278174551587662557388862052117599855872835584;
            6'd29: xpb[46] = 256'd9837804457449558062072379053218752395071287221934438464268264656993582579712;
            6'd30: xpb[46] = 256'd10177039093913335926281771434364226615590986781311488066484411714131292323840;
            6'd31: xpb[46] = 256'd10516273730377113790491163815509700836110686340688537668700558771269002067968;
            6'd32: xpb[46] = 256'd10855508366840891654700556196655175056630385900065587270916705828406711812096;
            6'd33: xpb[46] = 256'd11194743003304669518909948577800649277150085459442636873132852885544421556224;
            6'd34: xpb[46] = 256'd11533977639768447383119340958946123497669785018819686475348999942682131300352;
            6'd35: xpb[46] = 256'd11873212276232225247328733340091597718189484578196736077565146999819841044480;
            6'd36: xpb[46] = 256'd12212446912696003111538125721237071938709184137573785679781294056957550788608;
            6'd37: xpb[46] = 256'd12551681549159780975747518102382546159228883696950835281997441114095260532736;
            6'd38: xpb[46] = 256'd12890916185623558839956910483528020379748583256327884884213588171232970276864;
            6'd39: xpb[46] = 256'd13230150822087336704166302864673494600268282815704934486429735228370680020992;
            6'd40: xpb[46] = 256'd13569385458551114568375695245818968820787982375081984088645882285508389765120;
            6'd41: xpb[46] = 256'd13908620095014892432585087626964443041307681934459033690862029342646099509248;
            6'd42: xpb[46] = 256'd14247854731478670296794480008109917261827381493836083293078176399783809253376;
            6'd43: xpb[46] = 256'd14587089367942448161003872389255391482347081053213132895294323456921518997504;
            6'd44: xpb[46] = 256'd14926324004406226025213264770400865702866780612590182497510470514059228741632;
            6'd45: xpb[46] = 256'd15265558640870003889422657151546339923386480171967232099726617571196938485760;
            6'd46: xpb[46] = 256'd15604793277333781753632049532691814143906179731344281701942764628334648229888;
            6'd47: xpb[46] = 256'd15944027913797559617841441913837288364425879290721331304158911685472357974016;
            6'd48: xpb[46] = 256'd16283262550261337482050834294982762584945578850098380906375058742610067718144;
            6'd49: xpb[46] = 256'd16622497186725115346260226676128236805465278409475430508591205799747777462272;
            6'd50: xpb[46] = 256'd16961731823188893210469619057273711025984977968852480110807352856885487206400;
            6'd51: xpb[46] = 256'd17300966459652671074679011438419185246504677528229529713023499914023196950528;
            6'd52: xpb[46] = 256'd17640201096116448938888403819564659467024377087606579315239646971160906694656;
            6'd53: xpb[46] = 256'd17979435732580226803097796200710133687544076646983628917455794028298616438784;
            6'd54: xpb[46] = 256'd18318670369044004667307188581855607908063776206360678519671941085436326182912;
            6'd55: xpb[46] = 256'd18657905005507782531516580963001082128583475765737728121888088142574035927040;
            6'd56: xpb[46] = 256'd18997139641971560395725973344146556349103175325114777724104235199711745671168;
            6'd57: xpb[46] = 256'd19336374278435338259935365725292030569622874884491827326320382256849455415296;
            6'd58: xpb[46] = 256'd19675608914899116124144758106437504790142574443868876928536529313987165159424;
            6'd59: xpb[46] = 256'd20014843551362893988354150487582979010662274003245926530752676371124874903552;
            6'd60: xpb[46] = 256'd20354078187826671852563542868728453231181973562622976132968823428262584647680;
            6'd61: xpb[46] = 256'd20693312824290449716772935249873927451701673122000025735184970485400294391808;
            6'd62: xpb[46] = 256'd21032547460754227580982327631019401672221372681377075337401117542538004135936;
            6'd63: xpb[46] = 256'd21371782097218005445191720012164875892741072240754124939617264599675713880064;
        endcase
    end

    always_comb begin
        case(flag[47])
            6'd0: xpb[47] = 256'd0;
            6'd1: xpb[47] = 256'd21711016733681783309401112393310350113260771800131174541833411656813423624192;
            6'd2: xpb[47] = 256'd43422033467363566618802224786620700226521543600262349083666823313626847248384;
            6'd3: xpb[47] = 256'd65133050201045349928203337179931050339782315400393523625500234970440270872576;
            6'd4: xpb[47] = 256'd86844066934727133237604449573241400453043087200524698167333646627253694496768;
            6'd5: xpb[47] = 256'd108555083668408916547005561966551750566303859000655872709167058284067118120960;
            6'd6: xpb[47] = 256'd14474011191734451099986329145841207913314276808862855796579276007590856753153;
            6'd7: xpb[47] = 256'd36185027925416234409387441539151558026575048608994030338412687664404280377345;
            6'd8: xpb[47] = 256'd57896044659098017718788553932461908139835820409125204880246099321217704001537;
            6'd9: xpb[47] = 256'd79607061392779801028189666325772258253096592209256379422079510978031127625729;
            6'd10: xpb[47] = 256'd101318078126461584337590778719082608366357364009387553963912922634844551249921;
            6'd11: xpb[47] = 256'd7237005649787118890571545898372065713367781817594537051325140358368289882114;
            6'd12: xpb[47] = 256'd28948022383468902199972658291682415826628553617725711593158552015181713506306;
            6'd13: xpb[47] = 256'd50659039117150685509373770684992765939889325417856886134991963671995137130498;
            6'd14: xpb[47] = 256'd72370055850832468818774883078303116053150097217988060676825375328808560754690;
            6'd15: xpb[47] = 256'd94081072584514252128175995471613466166410869018119235218658786985621984378882;
            6'd16: xpb[47] = 256'd107839786681156762650902923513421286826326218306071004709145723011075;
            6'd17: xpb[47] = 256'd21711016841521569990557875044213273626682058626457392847904416365959146635267;
            6'd18: xpb[47] = 256'd43422033575203353299958987437523623739942830426588567389737828022772570259459;
            6'd19: xpb[47] = 256'd65133050308885136609360099830833973853203602226719741931571239679585993883651;
            6'd20: xpb[47] = 256'd86844067042566919918761212224144323966464374026850916473404651336399417507843;
            6'd21: xpb[47] = 256'd108555083776248703228162324617454674079725145826982091015238062993212841132035;
            6'd22: xpb[47] = 256'd14474011299574237781143091796744131426735563635189074102650280716736579764228;
            6'd23: xpb[47] = 256'd36185028033256021090544204190054481539996335435320248644483692373550003388420;
            6'd24: xpb[47] = 256'd57896044766937804399945316583364831653257107235451423186317104030363427012612;
            6'd25: xpb[47] = 256'd79607061500619587709346428976675181766517879035582597728150515687176850636804;
            6'd26: xpb[47] = 256'd101318078234301371018747541369985531879778650835713772269983927343990274260996;
            6'd27: xpb[47] = 256'd7237005757626905571728308549274989226789068643920755357396145067514012893189;
            6'd28: xpb[47] = 256'd28948022491308688881129420942585339340049840444051929899229556724327436517381;
            6'd29: xpb[47] = 256'd50659039224990472190530533335895689453310612244183104441062968381140860141573;
            6'd30: xpb[47] = 256'd72370055958672255499931645729206039566571384044314278982896380037954283765765;
            6'd31: xpb[47] = 256'd94081072692354038809332758122516389679832155844445453524729791694767707389957;
            6'd32: xpb[47] = 256'd215679573362313525301805847026842573652652436612142009418291446022150;
            6'd33: xpb[47] = 256'd21711016949361356671714637695116197140103345452783611153975421075104869646342;
            6'd34: xpb[47] = 256'd43422033683043139981115750088426547253364117252914785695808832731918293270534;
            6'd35: xpb[47] = 256'd65133050416724923290516862481736897366624889053045960237642244388731716894726;
            6'd36: xpb[47] = 256'd86844067150406706599917974875047247479885660853177134779475656045545140518918;
            6'd37: xpb[47] = 256'd108555083884088489909319087268357597593146432653308309321309067702358564143110;
            6'd38: xpb[47] = 256'd14474011407414024462299854447647054940156850461515292408721285425882302775303;
            6'd39: xpb[47] = 256'd36185028141095807771700966840957405053417622261646466950554697082695726399495;
            6'd40: xpb[47] = 256'd57896044874777591081102079234267755166678394061777641492388108739509150023687;
            6'd41: xpb[47] = 256'd79607061608459374390503191627578105279939165861908816034221520396322573647879;
            6'd42: xpb[47] = 256'd101318078342141157699904304020888455393199937662039990576054932053135997272071;
            6'd43: xpb[47] = 256'd7237005865466692252885071200177912740210355470246973663467149776659735904264;
            6'd44: xpb[47] = 256'd28948022599148475562286183593488262853471127270378148205300561433473159528456;
            6'd45: xpb[47] = 256'd50659039332830258871687295986798612966731899070509322747133973090286583152648;
            6'd46: xpb[47] = 256'd72370056066512042181088408380108963079992670870640497288967384747100006776840;
            6'd47: xpb[47] = 256'd94081072800193825490489520773419313193253442670771671830800796403913430401032;
            6'd48: xpb[47] = 256'd323519360043470287952708770540263860478978654918213014127437169033225;
            6'd49: xpb[47] = 256'd21711017057201143352871400346019120653524632279109829460046425784250592657417;
            6'd50: xpb[47] = 256'd43422033790882926662272512739329470766785404079241004001879837441064016281609;
            6'd51: xpb[47] = 256'd65133050524564709971673625132639820880046175879372178543713249097877439905801;
            6'd52: xpb[47] = 256'd86844067258246493281074737525950170993306947679503353085546660754690863529993;
            6'd53: xpb[47] = 256'd108555083991928276590475849919260521106567719479634527627380072411504287154185;
            6'd54: xpb[47] = 256'd14474011515253811143456617098549978453578137287841510714792290135028025786378;
            6'd55: xpb[47] = 256'd36185028248935594452857729491860328566838909087972685256625701791841449410570;
            6'd56: xpb[47] = 256'd57896044982617377762258841885170678680099680888103859798459113448654873034762;
            6'd57: xpb[47] = 256'd79607061716299161071659954278481028793360452688235034340292525105468296658954;
            6'd58: xpb[47] = 256'd101318078449980944381061066671791378906621224488366208882125936762281720283146;
            6'd59: xpb[47] = 256'd7237005973306478934041833851080836253631642296573191969538154485805458915339;
            6'd60: xpb[47] = 256'd28948022706988262243442946244391186366892414096704366511371566142618882539531;
            6'd61: xpb[47] = 256'd50659039440670045552844058637701536480153185896835541053204977799432306163723;
            6'd62: xpb[47] = 256'd72370056174351828862245171031011886593413957696966715595038389456245729787915;
            6'd63: xpb[47] = 256'd94081072908033612171646283424322236706674729497097890136871801113059153412107;
        endcase
    end

    always_comb begin
        case(flag[48])
            6'd0: xpb[48] = 256'd0;
            6'd1: xpb[48] = 256'd107839786681156762650902923513421286826326218306071004709145723011075;
            6'd2: xpb[48] = 256'd215679573362313525301805847026842573652652436612142009418291446022150;
            6'd3: xpb[48] = 256'd323519360043470287952708770540263860478978654918213014127437169033225;
            6'd4: xpb[48] = 256'd431359146724627050603611694053685147305304873224284018836582892044300;
            6'd5: xpb[48] = 256'd539198933405783813254514617567106434131631091530355023545728615055375;
            6'd6: xpb[48] = 256'd647038720086940575905417541080527720957957309836426028254874338066450;
            6'd7: xpb[48] = 256'd754878506768097338556320464593949007784283528142497032964020061077525;
            6'd8: xpb[48] = 256'd862718293449254101207223388107370294610609746448568037673165784088600;
            6'd9: xpb[48] = 256'd970558080130410863858126311620791581436935964754639042382311507099675;
            6'd10: xpb[48] = 256'd1078397866811567626509029235134212868263262183060710047091457230110750;
            6'd11: xpb[48] = 256'd1186237653492724389159932158647634155089588401366781051800602953121825;
            6'd12: xpb[48] = 256'd1294077440173881151810835082161055441915914619672852056509748676132900;
            6'd13: xpb[48] = 256'd1401917226855037914461738005674476728742240837978923061218894399143975;
            6'd14: xpb[48] = 256'd1509757013536194677112640929187898015568567056284994065928040122155050;
            6'd15: xpb[48] = 256'd1617596800217351439763543852701319302394893274591065070637185845166125;
            6'd16: xpb[48] = 256'd1725436586898508202414446776214740589221219492897136075346331568177200;
            6'd17: xpb[48] = 256'd1833276373579664965065349699728161876047545711203207080055477291188275;
            6'd18: xpb[48] = 256'd1941116160260821727716252623241583162873871929509278084764623014199350;
            6'd19: xpb[48] = 256'd2048955946941978490367155546755004449700198147815349089473768737210425;
            6'd20: xpb[48] = 256'd2156795733623135253018058470268425736526524366121420094182914460221500;
            6'd21: xpb[48] = 256'd2264635520304292015668961393781847023352850584427491098892060183232575;
            6'd22: xpb[48] = 256'd2372475306985448778319864317295268310179176802733562103601205906243650;
            6'd23: xpb[48] = 256'd2480315093666605540970767240808689597005503021039633108310351629254725;
            6'd24: xpb[48] = 256'd2588154880347762303621670164322110883831829239345704113019497352265800;
            6'd25: xpb[48] = 256'd2695994667028919066272573087835532170658155457651775117728643075276875;
            6'd26: xpb[48] = 256'd2803834453710075828923476011348953457484481675957846122437788798287950;
            6'd27: xpb[48] = 256'd2911674240391232591574378934862374744310807894263917127146934521299025;
            6'd28: xpb[48] = 256'd3019514027072389354225281858375796031137134112569988131856080244310100;
            6'd29: xpb[48] = 256'd3127353813753546116876184781889217317963460330876059136565225967321175;
            6'd30: xpb[48] = 256'd3235193600434702879527087705402638604789786549182130141274371690332250;
            6'd31: xpb[48] = 256'd3343033387115859642177990628916059891616112767488201145983517413343325;
            6'd32: xpb[48] = 256'd3450873173797016404828893552429481178442438985794272150692663136354400;
            6'd33: xpb[48] = 256'd3558712960478173167479796475942902465268765204100343155401808859365475;
            6'd34: xpb[48] = 256'd3666552747159329930130699399456323752095091422406414160110954582376550;
            6'd35: xpb[48] = 256'd3774392533840486692781602322969745038921417640712485164820100305387625;
            6'd36: xpb[48] = 256'd3882232320521643455432505246483166325747743859018556169529246028398700;
            6'd37: xpb[48] = 256'd3990072107202800218083408169996587612574070077324627174238391751409775;
            6'd38: xpb[48] = 256'd4097911893883956980734311093510008899400396295630698178947537474420850;
            6'd39: xpb[48] = 256'd4205751680565113743385214017023430186226722513936769183656683197431925;
            6'd40: xpb[48] = 256'd4313591467246270506036116940536851473053048732242840188365828920443000;
            6'd41: xpb[48] = 256'd4421431253927427268687019864050272759879374950548911193074974643454075;
            6'd42: xpb[48] = 256'd4529271040608584031337922787563694046705701168854982197784120366465150;
            6'd43: xpb[48] = 256'd4637110827289740793988825711077115333532027387161053202493266089476225;
            6'd44: xpb[48] = 256'd4744950613970897556639728634590536620358353605467124207202411812487300;
            6'd45: xpb[48] = 256'd4852790400652054319290631558103957907184679823773195211911557535498375;
            6'd46: xpb[48] = 256'd4960630187333211081941534481617379194011006042079266216620703258509450;
            6'd47: xpb[48] = 256'd5068469974014367844592437405130800480837332260385337221329848981520525;
            6'd48: xpb[48] = 256'd5176309760695524607243340328644221767663658478691408226038994704531600;
            6'd49: xpb[48] = 256'd5284149547376681369894243252157643054489984696997479230748140427542675;
            6'd50: xpb[48] = 256'd5391989334057838132545146175671064341316310915303550235457286150553750;
            6'd51: xpb[48] = 256'd5499829120738994895196049099184485628142637133609621240166431873564825;
            6'd52: xpb[48] = 256'd5607668907420151657846952022697906914968963351915692244875577596575900;
            6'd53: xpb[48] = 256'd5715508694101308420497854946211328201795289570221763249584723319586975;
            6'd54: xpb[48] = 256'd5823348480782465183148757869724749488621615788527834254293869042598050;
            6'd55: xpb[48] = 256'd5931188267463621945799660793238170775447942006833905259003014765609125;
            6'd56: xpb[48] = 256'd6039028054144778708450563716751592062274268225139976263712160488620200;
            6'd57: xpb[48] = 256'd6146867840825935471101466640265013349100594443446047268421306211631275;
            6'd58: xpb[48] = 256'd6254707627507092233752369563778434635926920661752118273130451934642350;
            6'd59: xpb[48] = 256'd6362547414188248996403272487291855922753246880058189277839597657653425;
            6'd60: xpb[48] = 256'd6470387200869405759054175410805277209579573098364260282548743380664500;
            6'd61: xpb[48] = 256'd6578226987550562521705078334318698496405899316670331287257889103675575;
            6'd62: xpb[48] = 256'd6686066774231719284355981257832119783232225534976402291967034826686650;
            6'd63: xpb[48] = 256'd6793906560912876047006884181345541070058551753282473296676180549697725;
        endcase
    end

    always_comb begin
        case(flag[49])
            6'd0: xpb[49] = 256'd0;
            6'd1: xpb[49] = 256'd6901746347594032809657787104858962356884877971588544301385326272708800;
            6'd2: xpb[49] = 256'd13803492695188065619315574209717924713769755943177088602770652545417600;
            6'd3: xpb[49] = 256'd20705239042782098428973361314576887070654633914765632904155978818126400;
            6'd4: xpb[49] = 256'd27606985390376131238631148419435849427539511886354177205541305090835200;
            6'd5: xpb[49] = 256'd34508731737970164048288935524294811784424389857942721506926631363544000;
            6'd6: xpb[49] = 256'd41410478085564196857946722629153774141309267829531265808311957636252800;
            6'd7: xpb[49] = 256'd48312224433158229667604509734012736498194145801119810109697283908961600;
            6'd8: xpb[49] = 256'd55213970780752262477262296838871698855079023772708354411082610181670400;
            6'd9: xpb[49] = 256'd62115717128346295286920083943730661211963901744296898712467936454379200;
            6'd10: xpb[49] = 256'd69017463475940328096577871048589623568848779715885443013853262727088000;
            6'd11: xpb[49] = 256'd75919209823534360906235658153448585925733657687473987315238588999796800;
            6'd12: xpb[49] = 256'd82820956171128393715893445258307548282618535659062531616623915272505600;
            6'd13: xpb[49] = 256'd89722702518722426525551232363166510639503413630651075918009241545214400;
            6'd14: xpb[49] = 256'd96624448866316459335209019468025472996388291602239620219394567817923200;
            6'd15: xpb[49] = 256'd103526195213910492144866806572884435353273169573828164520779894090632000;
            6'd16: xpb[49] = 256'd110427941561504524954524593677743397710158047545416708822165220363340800;
            6'd17: xpb[49] = 256'd117329687909098557764182380782602360067042925517005253123550546636049600;
            6'd18: xpb[49] = 256'd124231434256692590573840167887461322423927803488593797424935872908758400;
            6'd19: xpb[49] = 256'd131133180604286623383497954992320284780812681460182341726321199181467200;
            6'd20: xpb[49] = 256'd138034926951880656193155742097179247137697559431770886027706525454176000;
            6'd21: xpb[49] = 256'd144936673299474689002813529202038209494582437403359430329091851726884800;
            6'd22: xpb[49] = 256'd151838419647068721812471316306897171851467315374947974630477177999593600;
            6'd23: xpb[49] = 256'd158740165994662754622129103411756134208352193346536518931862504272302400;
            6'd24: xpb[49] = 256'd165641912342256787431786890516615096565237071318125063233247830545011200;
            6'd25: xpb[49] = 256'd172543658689850820241444677621474058922121949289713607534633156817720000;
            6'd26: xpb[49] = 256'd179445405037444853051102464726333021279006827261302151836018483090428800;
            6'd27: xpb[49] = 256'd186347151385038885860760251831191983635891705232890696137403809363137600;
            6'd28: xpb[49] = 256'd193248897732632918670418038936050945992776583204479240438789135635846400;
            6'd29: xpb[49] = 256'd200150644080226951480075826040909908349661461176067784740174461908555200;
            6'd30: xpb[49] = 256'd207052390427820984289733613145768870706546339147656329041559788181264000;
            6'd31: xpb[49] = 256'd213954136775415017099391400250627833063431217119244873342945114453972800;
            6'd32: xpb[49] = 256'd220855883123009049909049187355486795420316095090833417644330440726681600;
            6'd33: xpb[49] = 256'd227757629470603082718706974460345757777200973062421961945715766999390400;
            6'd34: xpb[49] = 256'd234659375818197115528364761565204720134085851034010506247101093272099200;
            6'd35: xpb[49] = 256'd241561122165791148338022548670063682490970729005599050548486419544808000;
            6'd36: xpb[49] = 256'd248462868513385181147680335774922644847855606977187594849871745817516800;
            6'd37: xpb[49] = 256'd255364614860979213957338122879781607204740484948776139151257072090225600;
            6'd38: xpb[49] = 256'd262266361208573246766995909984640569561625362920364683452642398362934400;
            6'd39: xpb[49] = 256'd269168107556167279576653697089499531918510240891953227754027724635643200;
            6'd40: xpb[49] = 256'd276069853903761312386311484194358494275395118863541772055413050908352000;
            6'd41: xpb[49] = 256'd282971600251355345195969271299217456632279996835130316356798377181060800;
            6'd42: xpb[49] = 256'd289873346598949378005627058404076418989164874806718860658183703453769600;
            6'd43: xpb[49] = 256'd296775092946543410815284845508935381346049752778307404959569029726478400;
            6'd44: xpb[49] = 256'd303676839294137443624942632613794343702934630749895949260954355999187200;
            6'd45: xpb[49] = 256'd310578585641731476434600419718653306059819508721484493562339682271896000;
            6'd46: xpb[49] = 256'd317480331989325509244258206823512268416704386693073037863725008544604800;
            6'd47: xpb[49] = 256'd324382078336919542053915993928371230773589264664661582165110334817313600;
            6'd48: xpb[49] = 256'd331283824684513574863573781033230193130474142636250126466495661090022400;
            6'd49: xpb[49] = 256'd338185571032107607673231568138089155487359020607838670767880987362731200;
            6'd50: xpb[49] = 256'd345087317379701640482889355242948117844243898579427215069266313635440000;
            6'd51: xpb[49] = 256'd351989063727295673292547142347807080201128776551015759370651639908148800;
            6'd52: xpb[49] = 256'd358890810074889706102204929452666042558013654522604303672036966180857600;
            6'd53: xpb[49] = 256'd365792556422483738911862716557525004914898532494192847973422292453566400;
            6'd54: xpb[49] = 256'd372694302770077771721520503662383967271783410465781392274807618726275200;
            6'd55: xpb[49] = 256'd379596049117671804531178290767242929628668288437369936576192944998984000;
            6'd56: xpb[49] = 256'd386497795465265837340836077872101891985553166408958480877578271271692800;
            6'd57: xpb[49] = 256'd393399541812859870150493864976960854342438044380547025178963597544401600;
            6'd58: xpb[49] = 256'd400301288160453902960151652081819816699322922352135569480348923817110400;
            6'd59: xpb[49] = 256'd407203034508047935769809439186678779056207800323724113781734250089819200;
            6'd60: xpb[49] = 256'd414104780855641968579467226291537741413092678295312658083119576362528000;
            6'd61: xpb[49] = 256'd421006527203236001389125013396396703769977556266901202384504902635236800;
            6'd62: xpb[49] = 256'd427908273550830034198782800501255666126862434238489746685890228907945600;
            6'd63: xpb[49] = 256'd434810019898424067008440587606114628483747312210078290987275555180654400;
        endcase
    end

    always_comb begin
        case(flag[50])
            6'd0: xpb[50] = 256'd0;
            6'd1: xpb[50] = 256'd441711766246018099818098374710973590840632190181666835288660881453363200;
            6'd2: xpb[50] = 256'd883423532492036199636196749421947181681264380363333670577321762906726400;
            6'd3: xpb[50] = 256'd1325135298738054299454295124132920772521896570545000505865982644360089600;
            6'd4: xpb[50] = 256'd1766847064984072399272393498843894363362528760726667341154643525813452800;
            6'd5: xpb[50] = 256'd2208558831230090499090491873554867954203160950908334176443304407266816000;
            6'd6: xpb[50] = 256'd2650270597476108598908590248265841545043793141090001011731965288720179200;
            6'd7: xpb[50] = 256'd3091982363722126698726688622976815135884425331271667847020626170173542400;
            6'd8: xpb[50] = 256'd3533694129968144798544786997687788726725057521453334682309287051626905600;
            6'd9: xpb[50] = 256'd3975405896214162898362885372398762317565689711635001517597947933080268800;
            6'd10: xpb[50] = 256'd4417117662460180998180983747109735908406321901816668352886608814533632000;
            6'd11: xpb[50] = 256'd4858829428706199097999082121820709499246954091998335188175269695986995200;
            6'd12: xpb[50] = 256'd5300541194952217197817180496531683090087586282180002023463930577440358400;
            6'd13: xpb[50] = 256'd5742252961198235297635278871242656680928218472361668858752591458893721600;
            6'd14: xpb[50] = 256'd6183964727444253397453377245953630271768850662543335694041252340347084800;
            6'd15: xpb[50] = 256'd6625676493690271497271475620664603862609482852725002529329913221800448000;
            6'd16: xpb[50] = 256'd7067388259936289597089573995375577453450115042906669364618574103253811200;
            6'd17: xpb[50] = 256'd7509100026182307696907672370086551044290747233088336199907234984707174400;
            6'd18: xpb[50] = 256'd7950811792428325796725770744797524635131379423270003035195895866160537600;
            6'd19: xpb[50] = 256'd8392523558674343896543869119508498225972011613451669870484556747613900800;
            6'd20: xpb[50] = 256'd8834235324920361996361967494219471816812643803633336705773217629067264000;
            6'd21: xpb[50] = 256'd9275947091166380096180065868930445407653275993815003541061878510520627200;
            6'd22: xpb[50] = 256'd9717658857412398195998164243641418998493908183996670376350539391973990400;
            6'd23: xpb[50] = 256'd10159370623658416295816262618352392589334540374178337211639200273427353600;
            6'd24: xpb[50] = 256'd10601082389904434395634360993063366180175172564360004046927861154880716800;
            6'd25: xpb[50] = 256'd11042794156150452495452459367774339771015804754541670882216522036334080000;
            6'd26: xpb[50] = 256'd11484505922396470595270557742485313361856436944723337717505182917787443200;
            6'd27: xpb[50] = 256'd11926217688642488695088656117196286952697069134905004552793843799240806400;
            6'd28: xpb[50] = 256'd12367929454888506794906754491907260543537701325086671388082504680694169600;
            6'd29: xpb[50] = 256'd12809641221134524894724852866618234134378333515268338223371165562147532800;
            6'd30: xpb[50] = 256'd13251352987380542994542951241329207725218965705450005058659826443600896000;
            6'd31: xpb[50] = 256'd13693064753626561094361049616040181316059597895631671893948487325054259200;
            6'd32: xpb[50] = 256'd14134776519872579194179147990751154906900230085813338729237148206507622400;
            6'd33: xpb[50] = 256'd14576488286118597293997246365462128497740862275995005564525809087960985600;
            6'd34: xpb[50] = 256'd15018200052364615393815344740173102088581494466176672399814469969414348800;
            6'd35: xpb[50] = 256'd15459911818610633493633443114884075679422126656358339235103130850867712000;
            6'd36: xpb[50] = 256'd15901623584856651593451541489595049270262758846540006070391791732321075200;
            6'd37: xpb[50] = 256'd16343335351102669693269639864306022861103391036721672905680452613774438400;
            6'd38: xpb[50] = 256'd16785047117348687793087738239016996451944023226903339740969113495227801600;
            6'd39: xpb[50] = 256'd17226758883594705892905836613727970042784655417085006576257774376681164800;
            6'd40: xpb[50] = 256'd17668470649840723992723934988438943633625287607266673411546435258134528000;
            6'd41: xpb[50] = 256'd18110182416086742092542033363149917224465919797448340246835096139587891200;
            6'd42: xpb[50] = 256'd18551894182332760192360131737860890815306551987630007082123757021041254400;
            6'd43: xpb[50] = 256'd18993605948578778292178230112571864406147184177811673917412417902494617600;
            6'd44: xpb[50] = 256'd19435317714824796391996328487282837996987816367993340752701078783947980800;
            6'd45: xpb[50] = 256'd19877029481070814491814426861993811587828448558175007587989739665401344000;
            6'd46: xpb[50] = 256'd20318741247316832591632525236704785178669080748356674423278400546854707200;
            6'd47: xpb[50] = 256'd20760453013562850691450623611415758769509712938538341258567061428308070400;
            6'd48: xpb[50] = 256'd21202164779808868791268721986126732360350345128720008093855722309761433600;
            6'd49: xpb[50] = 256'd21643876546054886891086820360837705951190977318901674929144383191214796800;
            6'd50: xpb[50] = 256'd22085588312300904990904918735548679542031609509083341764433044072668160000;
            6'd51: xpb[50] = 256'd22527300078546923090723017110259653132872241699265008599721704954121523200;
            6'd52: xpb[50] = 256'd22969011844792941190541115484970626723712873889446675435010365835574886400;
            6'd53: xpb[50] = 256'd23410723611038959290359213859681600314553506079628342270299026717028249600;
            6'd54: xpb[50] = 256'd23852435377284977390177312234392573905394138269810009105587687598481612800;
            6'd55: xpb[50] = 256'd24294147143530995489995410609103547496234770459991675940876348479934976000;
            6'd56: xpb[50] = 256'd24735858909777013589813508983814521087075402650173342776165009361388339200;
            6'd57: xpb[50] = 256'd25177570676023031689631607358525494677916034840355009611453670242841702400;
            6'd58: xpb[50] = 256'd25619282442269049789449705733236468268756667030536676446742331124295065600;
            6'd59: xpb[50] = 256'd26060994208515067889267804107947441859597299220718343282030992005748428800;
            6'd60: xpb[50] = 256'd26502705974761085989085902482658415450437931410900010117319652887201792000;
            6'd61: xpb[50] = 256'd26944417741007104088904000857369389041278563601081676952608313768655155200;
            6'd62: xpb[50] = 256'd27386129507253122188722099232080362632119195791263343787896974650108518400;
            6'd63: xpb[50] = 256'd27827841273499140288540197606791336222959827981445010623185635531561881600;
        endcase
    end

    always_comb begin
        case(flag[51])
            6'd0: xpb[51] = 256'd0;
            6'd1: xpb[51] = 256'd7067388259936289597089573995375577453450115042906669364618574103253811200;
            6'd2: xpb[51] = 256'd14134776519872579194179147990751154906900230085813338729237148206507622400;
            6'd3: xpb[51] = 256'd21202164779808868791268721986126732360350345128720008093855722309761433600;
            6'd4: xpb[51] = 256'd28269553039745158388358295981502309813800460171626677458474296413015244800;
            6'd5: xpb[51] = 256'd35336941299681447985447869976877887267250575214533346823092870516269056000;
            6'd6: xpb[51] = 256'd42404329559617737582537443972253464720700690257440016187711444619522867200;
            6'd7: xpb[51] = 256'd49471717819554027179627017967629042174150805300346685552330018722776678400;
            6'd8: xpb[51] = 256'd56539106079490316776716591963004619627600920343253354916948592826030489600;
            6'd9: xpb[51] = 256'd63606494339426606373806165958380197081051035386160024281567166929284300800;
            6'd10: xpb[51] = 256'd70673882599362895970895739953755774534501150429066693646185741032538112000;
            6'd11: xpb[51] = 256'd77741270859299185567985313949131351987951265471973363010804315135791923200;
            6'd12: xpb[51] = 256'd84808659119235475165074887944506929441401380514880032375422889239045734400;
            6'd13: xpb[51] = 256'd91876047379171764762164461939882506894851495557786701740041463342299545600;
            6'd14: xpb[51] = 256'd98943435639108054359254035935258084348301610600693371104660037445553356800;
            6'd15: xpb[51] = 256'd106010823899044343956343609930633661801751725643600040469278611548807168000;
            6'd16: xpb[51] = 256'd113078212158980633553433183926009239255201840686506709833897185652060979200;
            6'd17: xpb[51] = 256'd120145600418916923150522757921384816708651955729413379198515759755314790400;
            6'd18: xpb[51] = 256'd127212988678853212747612331916760394162102070772320048563134333858568601600;
            6'd19: xpb[51] = 256'd134280376938789502344701905912135971615552185815226717927752907961822412800;
            6'd20: xpb[51] = 256'd141347765198725791941791479907511549069002300858133387292371482065076224000;
            6'd21: xpb[51] = 256'd148415153458662081538881053902887126522452415901040056656990056168330035200;
            6'd22: xpb[51] = 256'd155482541718598371135970627898262703975902530943946726021608630271583846400;
            6'd23: xpb[51] = 256'd162549929978534660733060201893638281429352645986853395386227204374837657600;
            6'd24: xpb[51] = 256'd169617318238470950330149775889013858882802761029760064750845778478091468800;
            6'd25: xpb[51] = 256'd176684706498407239927239349884389436336252876072666734115464352581345280000;
            6'd26: xpb[51] = 256'd183752094758343529524328923879765013789702991115573403480082926684599091200;
            6'd27: xpb[51] = 256'd190819483018279819121418497875140591243153106158480072844701500787852902400;
            6'd28: xpb[51] = 256'd197886871278216108718508071870516168696603221201386742209320074891106713600;
            6'd29: xpb[51] = 256'd204954259538152398315597645865891746150053336244293411573938648994360524800;
            6'd30: xpb[51] = 256'd212021647798088687912687219861267323603503451287200080938557223097614336000;
            6'd31: xpb[51] = 256'd219089036058024977509776793856642901056953566330106750303175797200868147200;
            6'd32: xpb[51] = 256'd226156424317961267106866367852018478510403681373013419667794371304121958400;
            6'd33: xpb[51] = 256'd233223812577897556703955941847394055963853796415920089032412945407375769600;
            6'd34: xpb[51] = 256'd240291200837833846301045515842769633417303911458826758397031519510629580800;
            6'd35: xpb[51] = 256'd247358589097770135898135089838145210870754026501733427761650093613883392000;
            6'd36: xpb[51] = 256'd254425977357706425495224663833520788324204141544640097126268667717137203200;
            6'd37: xpb[51] = 256'd261493365617642715092314237828896365777654256587546766490887241820391014400;
            6'd38: xpb[51] = 256'd268560753877579004689403811824271943231104371630453435855505815923644825600;
            6'd39: xpb[51] = 256'd275628142137515294286493385819647520684554486673360105220124390026898636800;
            6'd40: xpb[51] = 256'd282695530397451583883582959815023098138004601716266774584742964130152448000;
            6'd41: xpb[51] = 256'd289762918657387873480672533810398675591454716759173443949361538233406259200;
            6'd42: xpb[51] = 256'd296830306917324163077762107805774253044904831802080113313980112336660070400;
            6'd43: xpb[51] = 256'd303897695177260452674851681801149830498354946844986782678598686439913881600;
            6'd44: xpb[51] = 256'd310965083437196742271941255796525407951805061887893452043217260543167692800;
            6'd45: xpb[51] = 256'd318032471697133031869030829791900985405255176930800121407835834646421504000;
            6'd46: xpb[51] = 256'd325099859957069321466120403787276562858705291973706790772454408749675315200;
            6'd47: xpb[51] = 256'd332167248217005611063209977782652140312155407016613460137072982852929126400;
            6'd48: xpb[51] = 256'd339234636476941900660299551778027717765605522059520129501691556956182937600;
            6'd49: xpb[51] = 256'd346302024736878190257389125773403295219055637102426798866310131059436748800;
            6'd50: xpb[51] = 256'd353369412996814479854478699768778872672505752145333468230928705162690560000;
            6'd51: xpb[51] = 256'd360436801256750769451568273764154450125955867188240137595547279265944371200;
            6'd52: xpb[51] = 256'd367504189516687059048657847759530027579405982231146806960165853369198182400;
            6'd53: xpb[51] = 256'd374571577776623348645747421754905605032856097274053476324784427472451993600;
            6'd54: xpb[51] = 256'd381638966036559638242836995750281182486306212316960145689403001575705804800;
            6'd55: xpb[51] = 256'd388706354296495927839926569745656759939756327359866815054021575678959616000;
            6'd56: xpb[51] = 256'd395773742556432217437016143741032337393206442402773484418640149782213427200;
            6'd57: xpb[51] = 256'd402841130816368507034105717736407914846656557445680153783258723885467238400;
            6'd58: xpb[51] = 256'd409908519076304796631195291731783492300106672488586823147877297988721049600;
            6'd59: xpb[51] = 256'd416975907336241086228284865727159069753556787531493492512495872091974860800;
            6'd60: xpb[51] = 256'd424043295596177375825374439722534647207006902574400161877114446195228672000;
            6'd61: xpb[51] = 256'd431110683856113665422464013717910224660457017617306831241733020298482483200;
            6'd62: xpb[51] = 256'd438178072116049955019553587713285802113907132660213500606351594401736294400;
            6'd63: xpb[51] = 256'd445245460375986244616643161708661379567357247703120169970970168504990105600;
        endcase
    end

    always_comb begin
        case(flag[52])
            6'd0: xpb[52] = 256'd0;
            6'd1: xpb[52] = 256'd452312848635922534213732735704036957020807362746026839335588742608243916800;
            6'd2: xpb[52] = 256'd904625697271845068427465471408073914041614725492053678671177485216487833600;
            6'd3: xpb[52] = 256'd1356938545907767602641198207112110871062422088238080518006766227824731750400;
            6'd4: xpb[52] = 256'd1809251394543690136854930942816147828083229450984107357342354970432975667200;
            6'd5: xpb[52] = 256'd2261564243179612671068663678520184785104036813730134196677943713041219584000;
            6'd6: xpb[52] = 256'd2713877091815535205282396414224221742124844176476161036013532455649463500800;
            6'd7: xpb[52] = 256'd3166189940451457739496129149928258699145651539222187875349121198257707417600;
            6'd8: xpb[52] = 256'd3618502789087380273709861885632295656166458901968214714684709940865951334400;
            6'd9: xpb[52] = 256'd4070815637723302807923594621336332613187266264714241554020298683474195251200;
            6'd10: xpb[52] = 256'd4523128486359225342137327357040369570208073627460268393355887426082439168000;
            6'd11: xpb[52] = 256'd4975441334995147876351060092744406527228880990206295232691476168690683084800;
            6'd12: xpb[52] = 256'd5427754183631070410564792828448443484249688352952322072027064911298927001600;
            6'd13: xpb[52] = 256'd5880067032266992944778525564152480441270495715698348911362653653907170918400;
            6'd14: xpb[52] = 256'd6332379880902915478992258299856517398291303078444375750698242396515414835200;
            6'd15: xpb[52] = 256'd6784692729538838013205991035560554355312110441190402590033831139123658752000;
            6'd16: xpb[52] = 256'd7237005578174760547419723771264591312332917803936429429369419881731902668800;
            6'd17: xpb[52] = 256'd7689318426810683081633456506968628269353725166682456268705008624340146585600;
            6'd18: xpb[52] = 256'd8141631275446605615847189242672665226374532529428483108040597366948390502400;
            6'd19: xpb[52] = 256'd8593944124082528150060921978376702183395339892174509947376186109556634419200;
            6'd20: xpb[52] = 256'd9046256972718450684274654714080739140416147254920536786711774852164878336000;
            6'd21: xpb[52] = 256'd9498569821354373218488387449784776097436954617666563626047363594773122252800;
            6'd22: xpb[52] = 256'd9950882669990295752702120185488813054457761980412590465382952337381366169600;
            6'd23: xpb[52] = 256'd10403195518626218286915852921192850011478569343158617304718541079989610086400;
            6'd24: xpb[52] = 256'd10855508367262140821129585656896886968499376705904644144054129822597854003200;
            6'd25: xpb[52] = 256'd11307821215898063355343318392600923925520184068650670983389718565206097920000;
            6'd26: xpb[52] = 256'd11760134064533985889557051128304960882540991431396697822725307307814341836800;
            6'd27: xpb[52] = 256'd12212446913169908423770783864008997839561798794142724662060896050422585753600;
            6'd28: xpb[52] = 256'd12664759761805830957984516599713034796582606156888751501396484793030829670400;
            6'd29: xpb[52] = 256'd13117072610441753492198249335417071753603413519634778340732073535639073587200;
            6'd30: xpb[52] = 256'd13569385459077676026411982071121108710624220882380805180067662278247317504000;
            6'd31: xpb[52] = 256'd14021698307713598560625714806825145667645028245126832019403251020855561420800;
            6'd32: xpb[52] = 256'd14474011156349521094839447542529182624665835607872858858738839763463805337600;
            6'd33: xpb[52] = 256'd14926324004985443629053180278233219581686642970618885698074428506072049254400;
            6'd34: xpb[52] = 256'd15378636853621366163266913013937256538707450333364912537410017248680293171200;
            6'd35: xpb[52] = 256'd15830949702257288697480645749641293495728257696110939376745605991288537088000;
            6'd36: xpb[52] = 256'd16283262550893211231694378485345330452749065058856966216081194733896781004800;
            6'd37: xpb[52] = 256'd16735575399529133765908111221049367409769872421602993055416783476505024921600;
            6'd38: xpb[52] = 256'd17187888248165056300121843956753404366790679784349019894752372219113268838400;
            6'd39: xpb[52] = 256'd17640201096800978834335576692457441323811487147095046734087960961721512755200;
            6'd40: xpb[52] = 256'd18092513945436901368549309428161478280832294509841073573423549704329756672000;
            6'd41: xpb[52] = 256'd18544826794072823902763042163865515237853101872587100412759138446938000588800;
            6'd42: xpb[52] = 256'd18997139642708746436976774899569552194873909235333127252094727189546244505600;
            6'd43: xpb[52] = 256'd19449452491344668971190507635273589151894716598079154091430315932154488422400;
            6'd44: xpb[52] = 256'd19901765339980591505404240370977626108915523960825180930765904674762732339200;
            6'd45: xpb[52] = 256'd20354078188616514039617973106681663065936331323571207770101493417370976256000;
            6'd46: xpb[52] = 256'd20806391037252436573831705842385700022957138686317234609437082159979220172800;
            6'd47: xpb[52] = 256'd21258703885888359108045438578089736979977946049063261448772670902587464089600;
            6'd48: xpb[52] = 256'd21711016734524281642259171313793773936998753411809288288108259645195708006400;
            6'd49: xpb[52] = 256'd22163329583160204176472904049497810894019560774555315127443848387803951923200;
            6'd50: xpb[52] = 256'd22615642431796126710686636785201847851040368137301341966779437130412195840000;
            6'd51: xpb[52] = 256'd23067955280432049244900369520905884808061175500047368806115025873020439756800;
            6'd52: xpb[52] = 256'd23520268129067971779114102256609921765081982862793395645450614615628683673600;
            6'd53: xpb[52] = 256'd23972580977703894313327834992313958722102790225539422484786203358236927590400;
            6'd54: xpb[52] = 256'd24424893826339816847541567728017995679123597588285449324121792100845171507200;
            6'd55: xpb[52] = 256'd24877206674975739381755300463722032636144404951031476163457380843453415424000;
            6'd56: xpb[52] = 256'd25329519523611661915969033199426069593165212313777503002792969586061659340800;
            6'd57: xpb[52] = 256'd25781832372247584450182765935130106550186019676523529842128558328669903257600;
            6'd58: xpb[52] = 256'd26234145220883506984396498670834143507206827039269556681464147071278147174400;
            6'd59: xpb[52] = 256'd26686458069519429518610231406538180464227634402015583520799735813886391091200;
            6'd60: xpb[52] = 256'd27138770918155352052823964142242217421248441764761610360135324556494635008000;
            6'd61: xpb[52] = 256'd27591083766791274587037696877946254378269249127507637199470913299102878924800;
            6'd62: xpb[52] = 256'd28043396615427197121251429613650291335290056490253664038806502041711122841600;
            6'd63: xpb[52] = 256'd28495709464063119655465162349354328292310863852999690878142090784319366758400;
        endcase
    end

    always_comb begin
        case(flag[53])
            6'd0: xpb[53] = 256'd0;
            6'd1: xpb[53] = 256'd28948022312699042189678895085058365249331671215745717717477679526927610675200;
            6'd2: xpb[53] = 256'd57896044625398084379357790170116730498663342431491435434955359053855221350400;
            6'd3: xpb[53] = 256'd86844066938097126569036685255175095747995013647237153152433038580782832025600;
            6'd4: xpb[53] = 256'd40439920002295235126212568231076330871058679415489524174420757708801;
            6'd5: xpb[53] = 256'd28948022353138962191974130211270933480408002086804397132967203701348368384001;
            6'd6: xpb[53] = 256'd57896044665838004381653025296329298729739673302550114850444883228275979059201;
            6'd7: xpb[53] = 256'd86844066978537046571331920381387663979071344518295832567922562755203589734401;
            6'd8: xpb[53] = 256'd80879840004590470252425136462152661742117358830979048348841515417602;
            6'd9: xpb[53] = 256'd28948022393578882194269365337483501711484332957863076548456727875769126092802;
            6'd10: xpb[53] = 256'd57896044706277924383948260422541866960816004173608794265934407402696736768002;
            6'd11: xpb[53] = 256'd86844067018976966573627155507600232210147675389354511983412086929624347443202;
            6'd12: xpb[53] = 256'd121319760006885705378637704693228992613176038246468572523262273126403;
            6'd13: xpb[53] = 256'd28948022434018802196564600463696069942560663828921755963946252050189883801603;
            6'd14: xpb[53] = 256'd57896044746717844386243495548754435191892335044667473681423931577117494476803;
            6'd15: xpb[53] = 256'd86844067059416886575922390633812800441224006260413191398901611104045105152003;
            6'd16: xpb[53] = 256'd161759680009180940504850272924305323484234717661958096697683030835204;
            6'd17: xpb[53] = 256'd28948022474458722198859835589908638173636994699980435379435776224610641510404;
            6'd18: xpb[53] = 256'd57896044787157764388538730674967003422968665915726153096913455751538252185604;
            6'd19: xpb[53] = 256'd86844067099856806578217625760025368672300337131471870814391135278465862860804;
            6'd20: xpb[53] = 256'd202199600011476175631062841155381654355293397077447620872103788544005;
            6'd21: xpb[53] = 256'd28948022514898642201155070716121206404713325571039114794925300399031399219205;
            6'd22: xpb[53] = 256'd57896044827597684390833965801179571654044996786784832512402979925959009894405;
            6'd23: xpb[53] = 256'd86844067140296726580512860886237936903376668002530550229880659452886620569605;
            6'd24: xpb[53] = 256'd242639520013771410757275409386457985226352076492937145046524546252806;
            6'd25: xpb[53] = 256'd28948022555338562203450305842333774635789656442097794210414824573452156928006;
            6'd26: xpb[53] = 256'd57896044868037604393129200927392139885121327657843511927892504100379767603206;
            6'd27: xpb[53] = 256'd86844067180736646582808096012450505134452998873589229645370183627307378278406;
            6'd28: xpb[53] = 256'd283079440016066645883487977617534316097410755908426669220945303961607;
            6'd29: xpb[53] = 256'd28948022595778482205745540968546342866865987313156473625904348747872914636807;
            6'd30: xpb[53] = 256'd57896044908477524395424436053604708116197658528902191343382028274800525312007;
            6'd31: xpb[53] = 256'd86844067221176566585103331138663073365529329744647909060859707801728135987207;
            6'd32: xpb[53] = 256'd323519360018361881009700545848610646968469435323916193395366061670408;
            6'd33: xpb[53] = 256'd28948022636218402208040776094758911097942318184215153041393872922293672345608;
            6'd34: xpb[53] = 256'd57896044948917444397719671179817276347273989399960870758871552449221283020808;
            6'd35: xpb[53] = 256'd86844067261616486587398566264875641596605660615706588476349231976148893696008;
            6'd36: xpb[53] = 256'd363959280020657116135913114079686977839528114739405717569786819379209;
            6'd37: xpb[53] = 256'd28948022676658322210336011220971479329018649055273832456883397096714430054409;
            6'd38: xpb[53] = 256'd57896044989357364400014906306029844578350320271019550174361076623642040729609;
            6'd39: xpb[53] = 256'd86844067302056406589693801391088209827681991486765267891838756150569651404809;
            6'd40: xpb[53] = 256'd404399200022952351262125682310763308710586794154895241744207577088010;
            6'd41: xpb[53] = 256'd28948022717098242212631246347184047560094979926332511872372921271135187763210;
            6'd42: xpb[53] = 256'd57896045029797284402310141432242412809426651142078229589850600798062798438410;
            6'd43: xpb[53] = 256'd86844067342496326591989036517300778058758322357823947307328280324990409113610;
            6'd44: xpb[53] = 256'd444839120025247586388338250541839639581645473570384765918628334796811;
            6'd45: xpb[53] = 256'd28948022757538162214926481473396615791171310797391191287862445445555945472011;
            6'd46: xpb[53] = 256'd57896045070237204404605376558454981040502982013136909005340124972483556147211;
            6'd47: xpb[53] = 256'd86844067382936246594284271643513346289834653228882626722817804499411166822411;
            6'd48: xpb[53] = 256'd485279040027542821514550818772915970452704152985874290093049092505612;
            6'd49: xpb[53] = 256'd28948022797978082217221716599609184022247641668449870703351969619976703180812;
            6'd50: xpb[53] = 256'd57896045110677124406900611684667549271579312884195588420829649146904313856012;
            6'd51: xpb[53] = 256'd86844067423376166596579506769725914520910984099941306138307328673831924531212;
            6'd52: xpb[53] = 256'd525718960029838056640763387003992301323762832401363814267469850214413;
            6'd53: xpb[53] = 256'd28948022838418002219516951725821752253323972539508550118841493794397460889613;
            6'd54: xpb[53] = 256'd57896045151117044409195846810880117502655643755254267836319173321325071564813;
            6'd55: xpb[53] = 256'd86844067463816086598874741895938482751987314970999985553796852848252682240013;
            6'd56: xpb[53] = 256'd566158880032133291766975955235068632194821511816853338441890607923214;
            6'd57: xpb[53] = 256'd28948022878857922221812186852034320484400303410567229534331017968818218598414;
            6'd58: xpb[53] = 256'd57896045191556964411491081937092685733731974626312947251808697495745829273614;
            6'd59: xpb[53] = 256'd86844067504256006601169977022151050983063645842058664969286377022673439948814;
            6'd60: xpb[53] = 256'd606598800034428526893188523466144963065880191232342862616311365632015;
            6'd61: xpb[53] = 256'd28948022919297842224107421978246888715476634281625908949820542143238976307215;
            6'd62: xpb[53] = 256'd57896045231996884413786317063305253964808305497371626667298221670166586982415;
            6'd63: xpb[53] = 256'd86844067544695926603465212148363619214139976713117344384775901197094197657615;
        endcase
    end

    always_comb begin
        case(flag[54])
            6'd0: xpb[54] = 256'd0;
            6'd1: xpb[54] = 256'd161759680009180940504850272924305323484234717661958096697683030835204;
            6'd2: xpb[54] = 256'd323519360018361881009700545848610646968469435323916193395366061670408;
            6'd3: xpb[54] = 256'd485279040027542821514550818772915970452704152985874290093049092505612;
            6'd4: xpb[54] = 256'd647038720036723762019401091697221293936938870647832386790732123340816;
            6'd5: xpb[54] = 256'd808798400045904702524251364621526617421173588309790483488415154176020;
            6'd6: xpb[54] = 256'd970558080055085643029101637545831940905408305971748580186098185011224;
            6'd7: xpb[54] = 256'd1132317760064266583533951910470137264389643023633706676883781215846428;
            6'd8: xpb[54] = 256'd1294077440073447524038802183394442587873877741295664773581464246681632;
            6'd9: xpb[54] = 256'd1455837120082628464543652456318747911358112458957622870279147277516836;
            6'd10: xpb[54] = 256'd1617596800091809405048502729243053234842347176619580966976830308352040;
            6'd11: xpb[54] = 256'd1779356480100990345553353002167358558326581894281539063674513339187244;
            6'd12: xpb[54] = 256'd1941116160110171286058203275091663881810816611943497160372196370022448;
            6'd13: xpb[54] = 256'd2102875840119352226563053548015969205295051329605455257069879400857652;
            6'd14: xpb[54] = 256'd2264635520128533167067903820940274528779286047267413353767562431692856;
            6'd15: xpb[54] = 256'd2426395200137714107572754093864579852263520764929371450465245462528060;
            6'd16: xpb[54] = 256'd2588154880146895048077604366788885175747755482591329547162928493363264;
            6'd17: xpb[54] = 256'd2749914560156075988582454639713190499231990200253287643860611524198468;
            6'd18: xpb[54] = 256'd2911674240165256929087304912637495822716224917915245740558294555033672;
            6'd19: xpb[54] = 256'd3073433920174437869592155185561801146200459635577203837255977585868876;
            6'd20: xpb[54] = 256'd3235193600183618810097005458486106469684694353239161933953660616704080;
            6'd21: xpb[54] = 256'd3396953280192799750601855731410411793168929070901120030651343647539284;
            6'd22: xpb[54] = 256'd3558712960201980691106706004334717116653163788563078127349026678374488;
            6'd23: xpb[54] = 256'd3720472640211161631611556277259022440137398506225036224046709709209692;
            6'd24: xpb[54] = 256'd3882232320220342572116406550183327763621633223886994320744392740044896;
            6'd25: xpb[54] = 256'd4043992000229523512621256823107633087105867941548952417442075770880100;
            6'd26: xpb[54] = 256'd4205751680238704453126107096031938410590102659210910514139758801715304;
            6'd27: xpb[54] = 256'd4367511360247885393630957368956243734074337376872868610837441832550508;
            6'd28: xpb[54] = 256'd4529271040257066334135807641880549057558572094534826707535124863385712;
            6'd29: xpb[54] = 256'd4691030720266247274640657914804854381042806812196784804232807894220916;
            6'd30: xpb[54] = 256'd4852790400275428215145508187729159704527041529858742900930490925056120;
            6'd31: xpb[54] = 256'd5014550080284609155650358460653465028011276247520700997628173955891324;
            6'd32: xpb[54] = 256'd5176309760293790096155208733577770351495510965182659094325856986726528;
            6'd33: xpb[54] = 256'd5338069440302971036660059006502075674979745682844617191023540017561732;
            6'd34: xpb[54] = 256'd5499829120312151977164909279426380998463980400506575287721223048396936;
            6'd35: xpb[54] = 256'd5661588800321332917669759552350686321948215118168533384418906079232140;
            6'd36: xpb[54] = 256'd5823348480330513858174609825274991645432449835830491481116589110067344;
            6'd37: xpb[54] = 256'd5985108160339694798679460098199296968916684553492449577814272140902548;
            6'd38: xpb[54] = 256'd6146867840348875739184310371123602292400919271154407674511955171737752;
            6'd39: xpb[54] = 256'd6308627520358056679689160644047907615885153988816365771209638202572956;
            6'd40: xpb[54] = 256'd6470387200367237620194010916972212939369388706478323867907321233408160;
            6'd41: xpb[54] = 256'd6632146880376418560698861189896518262853623424140281964605004264243364;
            6'd42: xpb[54] = 256'd6793906560385599501203711462820823586337858141802240061302687295078568;
            6'd43: xpb[54] = 256'd6955666240394780441708561735745128909822092859464198158000370325913772;
            6'd44: xpb[54] = 256'd7117425920403961382213412008669434233306327577126156254698053356748976;
            6'd45: xpb[54] = 256'd7279185600413142322718262281593739556790562294788114351395736387584180;
            6'd46: xpb[54] = 256'd7440945280422323263223112554518044880274797012450072448093419418419384;
            6'd47: xpb[54] = 256'd7602704960431504203727962827442350203759031730112030544791102449254588;
            6'd48: xpb[54] = 256'd7764464640440685144232813100366655527243266447773988641488785480089792;
            6'd49: xpb[54] = 256'd7926224320449866084737663373290960850727501165435946738186468510924996;
            6'd50: xpb[54] = 256'd8087984000459047025242513646215266174211735883097904834884151541760200;
            6'd51: xpb[54] = 256'd8249743680468227965747363919139571497695970600759862931581834572595404;
            6'd52: xpb[54] = 256'd8411503360477408906252214192063876821180205318421821028279517603430608;
            6'd53: xpb[54] = 256'd8573263040486589846757064464988182144664440036083779124977200634265812;
            6'd54: xpb[54] = 256'd8735022720495770787261914737912487468148674753745737221674883665101016;
            6'd55: xpb[54] = 256'd8896782400504951727766765010836792791632909471407695318372566695936220;
            6'd56: xpb[54] = 256'd9058542080514132668271615283761098115117144189069653415070249726771424;
            6'd57: xpb[54] = 256'd9220301760523313608776465556685403438601378906731611511767932757606628;
            6'd58: xpb[54] = 256'd9382061440532494549281315829609708762085613624393569608465615788441832;
            6'd59: xpb[54] = 256'd9543821120541675489786166102534014085569848342055527705163298819277036;
            6'd60: xpb[54] = 256'd9705580800550856430291016375458319409054083059717485801860981850112240;
            6'd61: xpb[54] = 256'd9867340480560037370795866648382624732538317777379443898558664880947444;
            6'd62: xpb[54] = 256'd10029100160569218311300716921306930056022552495041401995256347911782648;
            6'd63: xpb[54] = 256'd10190859840578399251805567194231235379506787212703360091954030942617852;
        endcase
    end

    always_comb begin
        case(flag[55])
            6'd0: xpb[55] = 256'd0;
            6'd1: xpb[55] = 256'd10352619520587580192310417467155540702991021930365318188651713973453056;
            6'd2: xpb[55] = 256'd20705239041175160384620834934311081405982043860730636377303427946906112;
            6'd3: xpb[55] = 256'd31057858561762740576931252401466622108973065791095954565955141920359168;
            6'd4: xpb[55] = 256'd41410478082350320769241669868622162811964087721461272754606855893812224;
            6'd5: xpb[55] = 256'd51763097602937900961552087335777703514955109651826590943258569867265280;
            6'd6: xpb[55] = 256'd62115717123525481153862504802933244217946131582191909131910283840718336;
            6'd7: xpb[55] = 256'd72468336644113061346172922270088784920937153512557227320561997814171392;
            6'd8: xpb[55] = 256'd82820956164700641538483339737244325623928175442922545509213711787624448;
            6'd9: xpb[55] = 256'd93173575685288221730793757204399866326919197373287863697865425761077504;
            6'd10: xpb[55] = 256'd103526195205875801923104174671555407029910219303653181886517139734530560;
            6'd11: xpb[55] = 256'd113878814726463382115414592138710947732901241234018500075168853707983616;
            6'd12: xpb[55] = 256'd124231434247050962307725009605866488435892263164383818263820567681436672;
            6'd13: xpb[55] = 256'd134584053767638542500035427073022029138883285094749136452472281654889728;
            6'd14: xpb[55] = 256'd144936673288226122692345844540177569841874307025114454641123995628342784;
            6'd15: xpb[55] = 256'd155289292808813702884656262007333110544865328955479772829775709601795840;
            6'd16: xpb[55] = 256'd165641912329401283076966679474488651247856350885845091018427423575248896;
            6'd17: xpb[55] = 256'd175994531849988863269277096941644191950847372816210409207079137548701952;
            6'd18: xpb[55] = 256'd186347151370576443461587514408799732653838394746575727395730851522155008;
            6'd19: xpb[55] = 256'd196699770891164023653897931875955273356829416676941045584382565495608064;
            6'd20: xpb[55] = 256'd207052390411751603846208349343110814059820438607306363773034279469061120;
            6'd21: xpb[55] = 256'd217405009932339184038518766810266354762811460537671681961685993442514176;
            6'd22: xpb[55] = 256'd227757629452926764230829184277421895465802482468037000150337707415967232;
            6'd23: xpb[55] = 256'd238110248973514344423139601744577436168793504398402318338989421389420288;
            6'd24: xpb[55] = 256'd248462868494101924615450019211732976871784526328767636527641135362873344;
            6'd25: xpb[55] = 256'd258815488014689504807760436678888517574775548259132954716292849336326400;
            6'd26: xpb[55] = 256'd269168107535277085000070854146044058277766570189498272904944563309779456;
            6'd27: xpb[55] = 256'd279520727055864665192381271613199598980757592119863591093596277283232512;
            6'd28: xpb[55] = 256'd289873346576452245384691689080355139683748614050228909282247991256685568;
            6'd29: xpb[55] = 256'd300225966097039825577002106547510680386739635980594227470899705230138624;
            6'd30: xpb[55] = 256'd310578585617627405769312524014666221089730657910959545659551419203591680;
            6'd31: xpb[55] = 256'd320931205138214985961622941481821761792721679841324863848203133177044736;
            6'd32: xpb[55] = 256'd331283824658802566153933358948977302495712701771690182036854847150497792;
            6'd33: xpb[55] = 256'd341636444179390146346243776416132843198703723702055500225506561123950848;
            6'd34: xpb[55] = 256'd351989063699977726538554193883288383901694745632420818414158275097403904;
            6'd35: xpb[55] = 256'd362341683220565306730864611350443924604685767562786136602809989070856960;
            6'd36: xpb[55] = 256'd372694302741152886923175028817599465307676789493151454791461703044310016;
            6'd37: xpb[55] = 256'd383046922261740467115485446284755006010667811423516772980113417017763072;
            6'd38: xpb[55] = 256'd393399541782328047307795863751910546713658833353882091168765130991216128;
            6'd39: xpb[55] = 256'd403752161302915627500106281219066087416649855284247409357416844964669184;
            6'd40: xpb[55] = 256'd414104780823503207692416698686221628119640877214612727546068558938122240;
            6'd41: xpb[55] = 256'd424457400344090787884727116153377168822631899144978045734720272911575296;
            6'd42: xpb[55] = 256'd434810019864678368077037533620532709525622921075343363923371986885028352;
            6'd43: xpb[55] = 256'd445162639385265948269347951087688250228613943005708682112023700858481408;
            6'd44: xpb[55] = 256'd455515258905853528461658368554843790931604964936074000300675414831934464;
            6'd45: xpb[55] = 256'd465867878426441108653968786021999331634595986866439318489327128805387520;
            6'd46: xpb[55] = 256'd476220497947028688846279203489154872337587008796804636677978842778840576;
            6'd47: xpb[55] = 256'd486573117467616269038589620956310413040578030727169954866630556752293632;
            6'd48: xpb[55] = 256'd496925736988203849230900038423465953743569052657535273055282270725746688;
            6'd49: xpb[55] = 256'd507278356508791429423210455890621494446560074587900591243933984699199744;
            6'd50: xpb[55] = 256'd517630976029379009615520873357777035149551096518265909432585698672652800;
            6'd51: xpb[55] = 256'd527983595549966589807831290824932575852542118448631227621237412646105856;
            6'd52: xpb[55] = 256'd538336215070554170000141708292088116555533140378996545809889126619558912;
            6'd53: xpb[55] = 256'd548688834591141750192452125759243657258524162309361863998540840593011968;
            6'd54: xpb[55] = 256'd559041454111729330384762543226399197961515184239727182187192554566465024;
            6'd55: xpb[55] = 256'd569394073632316910577072960693554738664506206170092500375844268539918080;
            6'd56: xpb[55] = 256'd579746693152904490769383378160710279367497228100457818564495982513371136;
            6'd57: xpb[55] = 256'd590099312673492070961693795627865820070488250030823136753147696486824192;
            6'd58: xpb[55] = 256'd600451932194079651154004213095021360773479271961188454941799410460277248;
            6'd59: xpb[55] = 256'd610804551714667231346314630562176901476470293891553773130451124433730304;
            6'd60: xpb[55] = 256'd621157171235254811538625048029332442179461315821919091319102838407183360;
            6'd61: xpb[55] = 256'd631509790755842391730935465496487982882452337752284409507754552380636416;
            6'd62: xpb[55] = 256'd641862410276429971923245882963643523585443359682649727696406266354089472;
            6'd63: xpb[55] = 256'd652215029797017552115556300430799064288434381613015045885057980327542528;
        endcase
    end

    always_comb begin
        case(flag[56])
            6'd0: xpb[56] = 256'd0;
            6'd1: xpb[56] = 256'd662567649317605132307866717897954604991425403543380364073709694300995584;
            6'd2: xpb[56] = 256'd1325135298635210264615733435795909209982850807086760728147419388601991168;
            6'd3: xpb[56] = 256'd1987702947952815396923600153693863814974276210630141092221129082902986752;
            6'd4: xpb[56] = 256'd2650270597270420529231466871591818419965701614173521456294838777203982336;
            6'd5: xpb[56] = 256'd3312838246588025661539333589489773024957127017716901820368548471504977920;
            6'd6: xpb[56] = 256'd3975405895905630793847200307387727629948552421260282184442258165805973504;
            6'd7: xpb[56] = 256'd4637973545223235926155067025285682234939977824803662548515967860106969088;
            6'd8: xpb[56] = 256'd5300541194540841058462933743183636839931403228347042912589677554407964672;
            6'd9: xpb[56] = 256'd5963108843858446190770800461081591444922828631890423276663387248708960256;
            6'd10: xpb[56] = 256'd6625676493176051323078667178979546049914254035433803640737096943009955840;
            6'd11: xpb[56] = 256'd7288244142493656455386533896877500654905679438977184004810806637310951424;
            6'd12: xpb[56] = 256'd7950811791811261587694400614775455259897104842520564368884516331611947008;
            6'd13: xpb[56] = 256'd8613379441128866720002267332673409864888530246063944732958226025912942592;
            6'd14: xpb[56] = 256'd9275947090446471852310134050571364469879955649607325097031935720213938176;
            6'd15: xpb[56] = 256'd9938514739764076984618000768469319074871381053150705461105645414514933760;
            6'd16: xpb[56] = 256'd10601082389081682116925867486367273679862806456694085825179355108815929344;
            6'd17: xpb[56] = 256'd11263650038399287249233734204265228284854231860237466189253064803116924928;
            6'd18: xpb[56] = 256'd11926217687716892381541600922163182889845657263780846553326774497417920512;
            6'd19: xpb[56] = 256'd12588785337034497513849467640061137494837082667324226917400484191718916096;
            6'd20: xpb[56] = 256'd13251352986352102646157334357959092099828508070867607281474193886019911680;
            6'd21: xpb[56] = 256'd13913920635669707778465201075857046704819933474410987645547903580320907264;
            6'd22: xpb[56] = 256'd14576488284987312910773067793755001309811358877954368009621613274621902848;
            6'd23: xpb[56] = 256'd15239055934304918043080934511652955914802784281497748373695322968922898432;
            6'd24: xpb[56] = 256'd15901623583622523175388801229550910519794209685041128737769032663223894016;
            6'd25: xpb[56] = 256'd16564191232940128307696667947448865124785635088584509101842742357524889600;
            6'd26: xpb[56] = 256'd17226758882257733440004534665346819729777060492127889465916452051825885184;
            6'd27: xpb[56] = 256'd17889326531575338572312401383244774334768485895671269829990161746126880768;
            6'd28: xpb[56] = 256'd18551894180892943704620268101142728939759911299214650194063871440427876352;
            6'd29: xpb[56] = 256'd19214461830210548836928134819040683544751336702758030558137581134728871936;
            6'd30: xpb[56] = 256'd19877029479528153969236001536938638149742762106301410922211290829029867520;
            6'd31: xpb[56] = 256'd20539597128845759101543868254836592754734187509844791286285000523330863104;
            6'd32: xpb[56] = 256'd21202164778163364233851734972734547359725612913388171650358710217631858688;
            6'd33: xpb[56] = 256'd21864732427480969366159601690632501964717038316931552014432419911932854272;
            6'd34: xpb[56] = 256'd22527300076798574498467468408530456569708463720474932378506129606233849856;
            6'd35: xpb[56] = 256'd23189867726116179630775335126428411174699889124018312742579839300534845440;
            6'd36: xpb[56] = 256'd23852435375433784763083201844326365779691314527561693106653548994835841024;
            6'd37: xpb[56] = 256'd24515003024751389895391068562224320384682739931105073470727258689136836608;
            6'd38: xpb[56] = 256'd25177570674068995027698935280122274989674165334648453834800968383437832192;
            6'd39: xpb[56] = 256'd25840138323386600160006801998020229594665590738191834198874678077738827776;
            6'd40: xpb[56] = 256'd26502705972704205292314668715918184199657016141735214562948387772039823360;
            6'd41: xpb[56] = 256'd27165273622021810424622535433816138804648441545278594927022097466340818944;
            6'd42: xpb[56] = 256'd27827841271339415556930402151714093409639866948821975291095807160641814528;
            6'd43: xpb[56] = 256'd28490408920657020689238268869612048014631292352365355655169516854942810112;
            6'd44: xpb[56] = 256'd29152976569974625821546135587510002619622717755908736019243226549243805696;
            6'd45: xpb[56] = 256'd29815544219292230953854002305407957224614143159452116383316936243544801280;
            6'd46: xpb[56] = 256'd30478111868609836086161869023305911829605568562995496747390645937845796864;
            6'd47: xpb[56] = 256'd31140679517927441218469735741203866434596993966538877111464355632146792448;
            6'd48: xpb[56] = 256'd31803247167245046350777602459101821039588419370082257475538065326447788032;
            6'd49: xpb[56] = 256'd32465814816562651483085469176999775644579844773625637839611775020748783616;
            6'd50: xpb[56] = 256'd33128382465880256615393335894897730249571270177169018203685484715049779200;
            6'd51: xpb[56] = 256'd33790950115197861747701202612795684854562695580712398567759194409350774784;
            6'd52: xpb[56] = 256'd34453517764515466880009069330693639459554120984255778931832904103651770368;
            6'd53: xpb[56] = 256'd35116085413833072012316936048591594064545546387799159295906613797952765952;
            6'd54: xpb[56] = 256'd35778653063150677144624802766489548669536971791342539659980323492253761536;
            6'd55: xpb[56] = 256'd36441220712468282276932669484387503274528397194885920024054033186554757120;
            6'd56: xpb[56] = 256'd37103788361785887409240536202285457879519822598429300388127742880855752704;
            6'd57: xpb[56] = 256'd37766356011103492541548402920183412484511248001972680752201452575156748288;
            6'd58: xpb[56] = 256'd38428923660421097673856269638081367089502673405516061116275162269457743872;
            6'd59: xpb[56] = 256'd39091491309738702806164136355979321694494098809059441480348871963758739456;
            6'd60: xpb[56] = 256'd39754058959056307938472003073877276299485524212602821844422581658059735040;
            6'd61: xpb[56] = 256'd40416626608373913070779869791775230904476949616146202208496291352360730624;
            6'd62: xpb[56] = 256'd41079194257691518203087736509673185509468375019689582572570001046661726208;
            6'd63: xpb[56] = 256'd41741761907009123335395603227571140114459800423232962936643710740962721792;
        endcase
    end



endmodule



